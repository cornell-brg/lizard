//-----------------------------------------------------------------------------
// proc
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.proc {"MemMsg": "MemMsg: op: 1 ts: 2 ad: 64 da: 8", "interface": ""}
// PyMTL: verilator_xinit = zeros
module proc
(
  input  logic [   0:0] clk,
  output logic [   0:0] db_recv_call,
  input  logic [  63:0] db_recv_msg,
  input  logic [   0:0] db_recv_rdy,
  output logic [   0:0] db_send_call,
  output logic [  63:0] db_send_msg,
  input  logic [   0:0] db_send_rdy,
  output logic [   0:0] mb_recv_0_call,
  input  logic [  75:0] mb_recv_0_msg,
  input  logic [   0:0] mb_recv_0_rdy,
  output logic [   0:0] mb_send_0_call,
  output logic [ 135:0] mb_send_0_msg,
  input  logic [   0:0] mb_send_0_rdy,
  input  logic [   0:0] reset
);

  // rename temporaries
  logic   [   1:0] rename$register_branch_mask;
  logic   [   5:0] rename$get_dst_preg;
  logic   [   4:0] rename$kill_notify_msg;
  logic   [ 189:0] rename$in_peek_msg;
  logic   [   0:0] rename$clk;
  logic   [   5:0] rename$get_src_preg$000;
  logic   [   5:0] rename$get_src_preg$001;
  logic   [   0:0] rename$get_dst_rdy;
  logic   [   0:0] rename$in_peek_rdy;
  logic   [   0:0] rename$register_spec_idx;
  logic   [   0:0] rename$reset;
  logic   [   0:0] rename$register_success;
  logic   [   0:0] rename$take_call;
  logic   [   3:0] rename$register_seq;
  logic   [   4:0] rename$get_src_areg$000;
  logic   [   4:0] rename$get_src_areg$001;
  logic   [   4:0] rename$get_dst_areg;
  logic   [  63:0] rename$register_pc;
  logic   [   0:0] rename$register_serialize;
  logic   [   0:0] rename$register_speculative;
  logic   [   0:0] rename$get_dst_call;
  logic   [   0:0] rename$register_call;
  logic   [ 141:0] rename$peek_msg;
  logic   [   0:0] rename$in_take_call;
  logic   [   0:0] rename$peek_rdy;
  logic   [  63:0] rename$register_pc_succ;

  GS11LRenameStage20LRenameDropController_0x6f71125cae5ffc5 rename
  (
    .register_branch_mask ( rename$register_branch_mask ),
    .get_dst_preg         ( rename$get_dst_preg ),
    .kill_notify_msg      ( rename$kill_notify_msg ),
    .in_peek_msg          ( rename$in_peek_msg ),
    .clk                  ( rename$clk ),
    .get_src_preg$000     ( rename$get_src_preg$000 ),
    .get_src_preg$001     ( rename$get_src_preg$001 ),
    .get_dst_rdy          ( rename$get_dst_rdy ),
    .in_peek_rdy          ( rename$in_peek_rdy ),
    .register_spec_idx    ( rename$register_spec_idx ),
    .reset                ( rename$reset ),
    .register_success     ( rename$register_success ),
    .take_call            ( rename$take_call ),
    .register_seq         ( rename$register_seq ),
    .get_src_areg$000     ( rename$get_src_areg$000 ),
    .get_src_areg$001     ( rename$get_src_areg$001 ),
    .get_dst_areg         ( rename$get_dst_areg ),
    .register_pc          ( rename$register_pc ),
    .register_serialize   ( rename$register_serialize ),
    .register_speculative ( rename$register_speculative ),
    .get_dst_call         ( rename$get_dst_call ),
    .register_call        ( rename$register_call ),
    .peek_msg             ( rename$peek_msg ),
    .in_take_call         ( rename$in_take_call ),
    .peek_rdy             ( rename$peek_rdy ),
    .register_pc_succ     ( rename$register_pc_succ )
  );

  // dispatch temporaries
  logic   [   4:0] dispatch$kill_notify_msg;
  logic   [ 141:0] dispatch$in_peek_msg;
  logic   [   0:0] dispatch$clk;
  logic   [   0:0] dispatch$in_peek_rdy;
  logic   [  63:0] dispatch$read_value$000;
  logic   [  63:0] dispatch$read_value$001;
  logic   [   0:0] dispatch$reset;
  logic   [   0:0] dispatch$take_call;
  logic   [ 250:0] dispatch$peek_msg;
  logic   [   0:0] dispatch$in_take_call;
  logic   [   0:0] dispatch$peek_rdy;
  logic   [   5:0] dispatch$read_tag$000;
  logic   [   5:0] dispatch$read_tag$001;

  GS13LDispatchStage22LDispatchDropController_0x78e60f5988db2eb3 dispatch
  (
    .kill_notify_msg ( dispatch$kill_notify_msg ),
    .in_peek_msg     ( dispatch$in_peek_msg ),
    .clk             ( dispatch$clk ),
    .in_peek_rdy     ( dispatch$in_peek_rdy ),
    .read_value$000  ( dispatch$read_value$000 ),
    .read_value$001  ( dispatch$read_value$001 ),
    .reset           ( dispatch$reset ),
    .take_call       ( dispatch$take_call ),
    .peek_msg        ( dispatch$peek_msg ),
    .in_take_call    ( dispatch$in_take_call ),
    .peek_rdy        ( dispatch$peek_rdy ),
    .read_tag$000    ( dispatch$read_tag$000 ),
    .read_tag$001    ( dispatch$read_tag$001 )
  );

  // alu temporaries
  logic   [   4:0] alu$kill_notify_msg;
  logic   [ 250:0] alu$in_peek_msg;
  logic   [   0:0] alu$clk;
  logic   [   0:0] alu$in_peek_rdy;
  logic   [   0:0] alu$reset;
  logic   [   0:0] alu$take_call;
  logic   [ 145:0] alu$peek_msg;
  logic   [   0:0] alu$in_take_call;
  logic   [   0:0] alu$peek_rdy;

  GS8LALUStage17LALUDropController_0xc628584b4321be9 alu
  (
    .kill_notify_msg ( alu$kill_notify_msg ),
    .in_peek_msg     ( alu$in_peek_msg ),
    .clk             ( alu$clk ),
    .in_peek_rdy     ( alu$in_peek_rdy ),
    .reset           ( alu$reset ),
    .take_call       ( alu$take_call ),
    .peek_msg        ( alu$peek_msg ),
    .in_take_call    ( alu$in_take_call ),
    .peek_rdy        ( alu$peek_rdy )
  );

  // decode temporaries
  logic   [   0:0] decode$kill_notify_msg;
  logic   [ 161:0] decode$in_peek_msg;
  logic   [   0:0] decode$clk;
  logic   [   0:0] decode$in_peek_rdy;
  logic   [   0:0] decode$reset;
  logic   [   0:0] decode$take_call;
  logic   [ 189:0] decode$peek_msg;
  logic   [   0:0] decode$in_take_call;
  logic   [   0:0] decode$peek_rdy;

  GS11LDecodeStage28LDecodeRedirectDropController_0x15fcfedd688afdf9 decode
  (
    .kill_notify_msg ( decode$kill_notify_msg ),
    .in_peek_msg     ( decode$in_peek_msg ),
    .clk             ( decode$clk ),
    .in_peek_rdy     ( decode$in_peek_rdy ),
    .reset           ( decode$reset ),
    .take_call       ( decode$take_call ),
    .peek_msg        ( decode$peek_msg ),
    .in_take_call    ( decode$in_take_call ),
    .peek_rdy        ( decode$peek_rdy )
  );

  // branch temporaries
  logic   [   4:0] branch$kill_notify_msg;
  logic   [ 250:0] branch$in_peek_msg;
  logic   [   0:0] branch$clk;
  logic   [   0:0] branch$in_peek_rdy;
  logic   [   0:0] branch$reset;
  logic   [   0:0] branch$take_call;
  logic   [   0:0] branch$cflow_redirect_call;
  logic   [  63:0] branch$cflow_redirect_target;
  logic   [ 145:0] branch$peek_msg;
  logic   [   3:0] branch$cflow_redirect_seq;
  logic   [   0:0] branch$cflow_redirect_force;
  logic   [   0:0] branch$in_take_call;
  logic   [   0:0] branch$peek_rdy;
  logic   [   0:0] branch$cflow_redirect_spec_idx;

  GS11LBranchStage20LBranchDropController_0xc628584b4321be9 branch
  (
    .kill_notify_msg         ( branch$kill_notify_msg ),
    .in_peek_msg             ( branch$in_peek_msg ),
    .clk                     ( branch$clk ),
    .in_peek_rdy             ( branch$in_peek_rdy ),
    .reset                   ( branch$reset ),
    .take_call               ( branch$take_call ),
    .cflow_redirect_call     ( branch$cflow_redirect_call ),
    .cflow_redirect_target   ( branch$cflow_redirect_target ),
    .peek_msg                ( branch$peek_msg ),
    .cflow_redirect_seq      ( branch$cflow_redirect_seq ),
    .cflow_redirect_force    ( branch$cflow_redirect_force ),
    .in_take_call            ( branch$in_take_call ),
    .peek_rdy                ( branch$peek_rdy ),
    .cflow_redirect_spec_idx ( branch$cflow_redirect_spec_idx )
  );

  // csr_pipe temporaries
  logic   [   4:0] csr_pipe$kill_notify_msg;
  logic   [ 250:0] csr_pipe$in_peek_msg;
  logic   [   0:0] csr_pipe$csr_op_success;
  logic   [  63:0] csr_pipe$csr_op_old;
  logic   [   0:0] csr_pipe$clk;
  logic   [   0:0] csr_pipe$in_peek_rdy;
  logic   [   0:0] csr_pipe$reset;
  logic   [   0:0] csr_pipe$take_call;
  logic   [   1:0] csr_pipe$csr_op_op;
  logic   [   0:0] csr_pipe$csr_op_call;
  logic   [   0:0] csr_pipe$csr_op_rs1_is_x0;
  logic   [ 145:0] csr_pipe$peek_msg;
  logic   [   0:0] csr_pipe$in_take_call;
  logic   [  11:0] csr_pipe$csr_op_csr;
  logic   [   0:0] csr_pipe$peek_rdy;
  logic   [  63:0] csr_pipe$csr_op_value;

  GS8LCSRStage17LCSRDropController_0xc628584b4321be9 csr_pipe
  (
    .kill_notify_msg  ( csr_pipe$kill_notify_msg ),
    .in_peek_msg      ( csr_pipe$in_peek_msg ),
    .csr_op_success   ( csr_pipe$csr_op_success ),
    .csr_op_old       ( csr_pipe$csr_op_old ),
    .clk              ( csr_pipe$clk ),
    .in_peek_rdy      ( csr_pipe$in_peek_rdy ),
    .reset            ( csr_pipe$reset ),
    .take_call        ( csr_pipe$take_call ),
    .csr_op_op        ( csr_pipe$csr_op_op ),
    .csr_op_call      ( csr_pipe$csr_op_call ),
    .csr_op_rs1_is_x0 ( csr_pipe$csr_op_rs1_is_x0 ),
    .peek_msg         ( csr_pipe$peek_msg ),
    .in_take_call     ( csr_pipe$in_take_call ),
    .csr_op_csr       ( csr_pipe$csr_op_csr ),
    .peek_rdy         ( csr_pipe$peek_rdy ),
    .csr_op_value     ( csr_pipe$csr_op_value )
  );

  // redirect_notifier temporaries
  logic   [   0:0] redirect_notifier$clk;
  logic   [  63:0] redirect_notifier$check_redirect_target;
  logic   [   0:0] redirect_notifier$reset;
  logic   [   0:0] redirect_notifier$check_redirect_redirect;
  logic   [   0:0] redirect_notifier$kill_notify_msg;

  RedirectNotifier_0x76bce5ec03c6a79c redirect_notifier
  (
    .clk                     ( redirect_notifier$clk ),
    .check_redirect_target   ( redirect_notifier$check_redirect_target ),
    .reset                   ( redirect_notifier$reset ),
    .check_redirect_redirect ( redirect_notifier$check_redirect_redirect ),
    .kill_notify_msg         ( redirect_notifier$kill_notify_msg )
  );

  // issue temporaries
  logic   [ 141:0] issue$in_peek_msg;
  logic   [   0:0] issue$clk;
  logic   [   4:0] issue$kill_notify_msg;
  logic   [   0:0] issue$in_peek_rdy;
  logic   [   0:0] issue$reset;
  logic   [   0:0] issue$is_ready_ready$000;
  logic   [   0:0] issue$is_ready_ready$001;
  logic   [  63:0] issue$get_updated_mask;
  logic   [   0:0] issue$take_call;
  logic   [   5:0] issue$is_ready_tag$000;
  logic   [   5:0] issue$is_ready_tag$001;
  logic   [ 141:0] issue$peek_msg;
  logic   [   0:0] issue$in_take_call;
  logic   [   0:0] issue$peek_rdy;

  Issue_0x52678fcc1604a432 issue
  (
    .in_peek_msg        ( issue$in_peek_msg ),
    .clk                ( issue$clk ),
    .kill_notify_msg    ( issue$kill_notify_msg ),
    .in_peek_rdy        ( issue$in_peek_rdy ),
    .reset              ( issue$reset ),
    .is_ready_ready$000 ( issue$is_ready_ready$000 ),
    .is_ready_ready$001 ( issue$is_ready_ready$001 ),
    .get_updated_mask   ( issue$get_updated_mask ),
    .take_call          ( issue$take_call ),
    .is_ready_tag$000   ( issue$is_ready_tag$000 ),
    .is_ready_tag$001   ( issue$is_ready_tag$001 ),
    .peek_msg           ( issue$peek_msg ),
    .in_take_call       ( issue$in_take_call ),
    .peek_rdy           ( issue$peek_rdy )
  );

  // csr temporaries
  logic   [  63:0] csr$debug_recv_msg;
  logic   [   0:0] csr$debug_recv_rdy;
  logic   [  11:0] csr$op_csr;
  logic   [   0:0] csr$debug_send_rdy;
  logic   [   0:0] csr$clk;
  logic   [   1:0] csr$op_op;
  logic   [   0:0] csr$op_call;
  logic   [   0:0] csr$op_rs1_is_x0;
  logic   [  63:0] csr$op_value;
  logic   [   0:0] csr$reset;
  logic   [   0:0] csr$debug_send_call;
  logic   [  63:0] csr$debug_send_msg;
  logic   [   0:0] csr$op_success;
  logic   [   0:0] csr$debug_recv_call;
  logic   [  63:0] csr$op_old;

  CSRManager_0x68582ff11a9d1315 csr
  (
    .debug_recv_msg  ( csr$debug_recv_msg ),
    .debug_recv_rdy  ( csr$debug_recv_rdy ),
    .op_csr          ( csr$op_csr ),
    .debug_send_rdy  ( csr$debug_send_rdy ),
    .clk             ( csr$clk ),
    .op_op           ( csr$op_op ),
    .op_call         ( csr$op_call ),
    .op_rs1_is_x0    ( csr$op_rs1_is_x0 ),
    .op_value        ( csr$op_value ),
    .reset           ( csr$reset ),
    .debug_send_call ( csr$debug_send_call ),
    .debug_send_msg  ( csr$debug_send_msg ),
    .op_success      ( csr$op_success ),
    .debug_recv_call ( csr$debug_recv_call ),
    .op_old          ( csr$op_old )
  );

  // writeback temporaries
  logic   [   4:0] writeback$kill_notify_msg;
  logic   [ 145:0] writeback$in_peek_msg;
  logic   [   0:0] writeback$clk;
  logic   [   0:0] writeback$in_peek_rdy;
  logic   [   0:0] writeback$reset;
  logic   [   0:0] writeback$take_call;
  logic   [   0:0] writeback$dataflow_write_call;
  logic   [ 141:0] writeback$peek_msg;
  logic   [   5:0] writeback$dataflow_write_tag;
  logic   [   0:0] writeback$in_take_call;
  logic   [  63:0] writeback$dataflow_write_value;
  logic   [   0:0] writeback$peek_rdy;

  GS14LWritebackStage23LWritebackDropController_0x4a102c6dab533550 writeback
  (
    .kill_notify_msg      ( writeback$kill_notify_msg ),
    .in_peek_msg          ( writeback$in_peek_msg ),
    .clk                  ( writeback$clk ),
    .in_peek_rdy          ( writeback$in_peek_rdy ),
    .reset                ( writeback$reset ),
    .take_call            ( writeback$take_call ),
    .dataflow_write_call  ( writeback$dataflow_write_call ),
    .peek_msg             ( writeback$peek_msg ),
    .dataflow_write_tag   ( writeback$dataflow_write_tag ),
    .in_take_call         ( writeback$in_take_call ),
    .dataflow_write_value ( writeback$dataflow_write_value ),
    .peek_rdy             ( writeback$peek_rdy )
  );

  // pipe_selector temporaries
  logic   [ 250:0] pipe_selector$in_peek_msg;
  logic   [   0:0] pipe_selector$branch_take_call;
  logic   [   0:0] pipe_selector$alu_take_call;
  logic   [   0:0] pipe_selector$clk;
  logic   [   0:0] pipe_selector$in_peek_rdy;
  logic   [   0:0] pipe_selector$reset;
  logic   [   0:0] pipe_selector$csr_take_call;
  logic   [ 250:0] pipe_selector$alu_peek_msg;
  logic   [   0:0] pipe_selector$branch_peek_rdy;
  logic   [   0:0] pipe_selector$alu_peek_rdy;
  logic   [ 250:0] pipe_selector$branch_peek_msg;
  logic   [   0:0] pipe_selector$in_take_call;
  logic   [   0:0] pipe_selector$csr_peek_rdy;
  logic   [ 250:0] pipe_selector$csr_peek_msg;

  PipeSelector_0x7f9520fbc84f298e pipe_selector
  (
    .in_peek_msg      ( pipe_selector$in_peek_msg ),
    .branch_take_call ( pipe_selector$branch_take_call ),
    .alu_take_call    ( pipe_selector$alu_take_call ),
    .clk              ( pipe_selector$clk ),
    .in_peek_rdy      ( pipe_selector$in_peek_rdy ),
    .reset            ( pipe_selector$reset ),
    .csr_take_call    ( pipe_selector$csr_take_call ),
    .alu_peek_msg     ( pipe_selector$alu_peek_msg ),
    .branch_peek_rdy  ( pipe_selector$branch_peek_rdy ),
    .alu_peek_rdy     ( pipe_selector$alu_peek_rdy ),
    .branch_peek_msg  ( pipe_selector$branch_peek_msg ),
    .in_take_call     ( pipe_selector$in_take_call ),
    .csr_peek_rdy     ( pipe_selector$csr_peek_rdy ),
    .csr_peek_msg     ( pipe_selector$csr_peek_msg )
  );

  // dflow temporaries
  logic   [   0:0] dflow$snapshot_call;
  logic   [   5:0] dflow$is_ready_tag$000;
  logic   [   5:0] dflow$is_ready_tag$001;
  logic   [   4:0] dflow$get_src_areg$000;
  logic   [   4:0] dflow$get_src_areg$001;
  logic   [   0:0] dflow$commit_call$000;
  logic   [   4:0] dflow$get_dst_areg$000;
  logic   [   5:0] dflow$write_tag$000;
  logic   [   0:0] dflow$get_dst_call$000;
  logic   [   0:0] dflow$restore_call;
  logic   [   0:0] dflow$clk;
  logic   [   0:0] dflow$write_call$000;
  logic   [   0:0] dflow$restore_source_id;
  logic   [  63:0] dflow$write_value$000;
  logic   [   0:0] dflow$free_snapshot_id_;
  logic   [   0:0] dflow$rollback_call;
  logic   [   0:0] dflow$free_snapshot_call;
  logic   [   0:0] dflow$reset;
  logic   [   5:0] dflow$read_tag$000;
  logic   [   5:0] dflow$read_tag$001;
  logic   [   5:0] dflow$commit_tag$000;
  logic   [   0:0] dflow$snapshot_rdy;
  logic   [   0:0] dflow$snapshot_id_;
  logic   [   5:0] dflow$get_dst_preg$000;
  logic   [   5:0] dflow$get_src_preg$000;
  logic   [   5:0] dflow$get_src_preg$001;
  logic   [   0:0] dflow$get_dst_rdy$000;
  logic   [  63:0] dflow$read_value$000;
  logic   [  63:0] dflow$read_value$001;
  logic   [   0:0] dflow$is_ready_ready$000;
  logic   [   0:0] dflow$is_ready_ready$001;
  logic   [  63:0] dflow$get_updated_mask;

  DataFlowManager_0x54912d9190dab9c9 dflow
  (
    .snapshot_call      ( dflow$snapshot_call ),
    .is_ready_tag$000   ( dflow$is_ready_tag$000 ),
    .is_ready_tag$001   ( dflow$is_ready_tag$001 ),
    .get_src_areg$000   ( dflow$get_src_areg$000 ),
    .get_src_areg$001   ( dflow$get_src_areg$001 ),
    .commit_call$000    ( dflow$commit_call$000 ),
    .get_dst_areg$000   ( dflow$get_dst_areg$000 ),
    .write_tag$000      ( dflow$write_tag$000 ),
    .get_dst_call$000   ( dflow$get_dst_call$000 ),
    .restore_call       ( dflow$restore_call ),
    .clk                ( dflow$clk ),
    .write_call$000     ( dflow$write_call$000 ),
    .restore_source_id  ( dflow$restore_source_id ),
    .write_value$000    ( dflow$write_value$000 ),
    .free_snapshot_id_  ( dflow$free_snapshot_id_ ),
    .rollback_call      ( dflow$rollback_call ),
    .free_snapshot_call ( dflow$free_snapshot_call ),
    .reset              ( dflow$reset ),
    .read_tag$000       ( dflow$read_tag$000 ),
    .read_tag$001       ( dflow$read_tag$001 ),
    .commit_tag$000     ( dflow$commit_tag$000 ),
    .snapshot_rdy       ( dflow$snapshot_rdy ),
    .snapshot_id_       ( dflow$snapshot_id_ ),
    .get_dst_preg$000   ( dflow$get_dst_preg$000 ),
    .get_src_preg$000   ( dflow$get_src_preg$000 ),
    .get_src_preg$001   ( dflow$get_src_preg$001 ),
    .get_dst_rdy$000    ( dflow$get_dst_rdy$000 ),
    .read_value$000     ( dflow$read_value$000 ),
    .read_value$001     ( dflow$read_value$001 ),
    .is_ready_ready$000 ( dflow$is_ready_ready$000 ),
    .is_ready_ready$001 ( dflow$is_ready_ready$001 ),
    .get_updated_mask   ( dflow$get_updated_mask )
  );

  // kill_notifier temporaries
  logic   [   0:0] kill_notifier$clk;
  logic   [   4:0] kill_notifier$check_kill_kill;
  logic   [   0:0] kill_notifier$reset;
  logic   [   4:0] kill_notifier$kill_notify_msg;

  KillNotifier_0x40986fce6fe74c56 kill_notifier
  (
    .clk             ( kill_notifier$clk ),
    .check_kill_kill ( kill_notifier$check_kill_kill ),
    .reset           ( kill_notifier$reset ),
    .kill_notify_msg ( kill_notifier$kill_notify_msg )
  );

  // writeback_arbiter temporaries
  logic   [ 145:0] writeback_arbiter$alu_peek_msg;
  logic   [   0:0] writeback_arbiter$clk;
  logic   [   0:0] writeback_arbiter$branch_peek_rdy;
  logic   [   0:0] writeback_arbiter$alu_peek_rdy;
  logic   [ 145:0] writeback_arbiter$branch_peek_msg;
  logic   [   0:0] writeback_arbiter$reset;
  logic   [   0:0] writeback_arbiter$csr_peek_rdy;
  logic   [ 145:0] writeback_arbiter$csr_peek_msg;
  logic   [   0:0] writeback_arbiter$take_call;
  logic   [   0:0] writeback_arbiter$branch_take_call;
  logic   [   0:0] writeback_arbiter$alu_take_call;
  logic   [ 145:0] writeback_arbiter$peek_msg;
  logic   [   0:0] writeback_arbiter$peek_rdy;
  logic   [   0:0] writeback_arbiter$csr_take_call;

  PipelineArbiter_0x311a0425acf3e6db writeback_arbiter
  (
    .alu_peek_msg     ( writeback_arbiter$alu_peek_msg ),
    .clk              ( writeback_arbiter$clk ),
    .branch_peek_rdy  ( writeback_arbiter$branch_peek_rdy ),
    .alu_peek_rdy     ( writeback_arbiter$alu_peek_rdy ),
    .branch_peek_msg  ( writeback_arbiter$branch_peek_msg ),
    .reset            ( writeback_arbiter$reset ),
    .csr_peek_rdy     ( writeback_arbiter$csr_peek_rdy ),
    .csr_peek_msg     ( writeback_arbiter$csr_peek_msg ),
    .take_call        ( writeback_arbiter$take_call ),
    .branch_take_call ( writeback_arbiter$branch_take_call ),
    .alu_take_call    ( writeback_arbiter$alu_take_call ),
    .peek_msg         ( writeback_arbiter$peek_msg ),
    .peek_rdy         ( writeback_arbiter$peek_rdy ),
    .csr_take_call    ( writeback_arbiter$csr_take_call )
  );

  // cflow temporaries
  logic   [   0:0] cflow$commit_call;
  logic   [   3:0] cflow$redirect_seq;
  logic   [  63:0] cflow$redirect_target;
  logic   [   0:0] cflow$redirect_call;
  logic   [   0:0] cflow$redirect_spec_idx;
  logic   [  63:0] cflow$register_pc_succ;
  logic   [   0:0] cflow$register_call;
  logic   [   0:0] cflow$clk;
  logic   [  63:0] cflow$register_pc;
  logic   [   0:0] cflow$register_speculative;
  logic   [   0:0] cflow$redirect_force;
  logic   [   0:0] cflow$dflow_snapshot_id_;
  logic   [   0:0] cflow$reset;
  logic   [   1:0] cflow$commit_status;
  logic   [   0:0] cflow$register_serialize;
  logic   [   0:0] cflow$dflow_snapshot_rdy;
  logic   [   4:0] cflow$check_kill_kill;
  logic   [   0:0] cflow$dflow_free_snapshot_id_;
  logic   [   0:0] cflow$dflow_restore_source_id;
  logic   [   3:0] cflow$get_head_seq;
  logic   [   0:0] cflow$register_success;
  logic   [   0:0] cflow$dflow_rollback_call;
  logic   [   0:0] cflow$dflow_snapshot_call;
  logic   [   0:0] cflow$register_spec_idx;
  logic   [  63:0] cflow$check_redirect_target;
  logic   [   0:0] cflow$dflow_free_snapshot_call;
  logic   [   0:0] cflow$check_redirect_redirect;
  logic   [   0:0] cflow$get_head_rdy;
  logic   [   1:0] cflow$register_branch_mask;
  logic   [   0:0] cflow$dflow_restore_call;
  logic   [   3:0] cflow$register_seq;

  ControlFlowManager_0x734ebf4161405225 cflow
  (
    .commit_call              ( cflow$commit_call ),
    .redirect_seq             ( cflow$redirect_seq ),
    .redirect_target          ( cflow$redirect_target ),
    .redirect_call            ( cflow$redirect_call ),
    .redirect_spec_idx        ( cflow$redirect_spec_idx ),
    .register_pc_succ         ( cflow$register_pc_succ ),
    .register_call            ( cflow$register_call ),
    .clk                      ( cflow$clk ),
    .register_pc              ( cflow$register_pc ),
    .register_speculative     ( cflow$register_speculative ),
    .redirect_force           ( cflow$redirect_force ),
    .dflow_snapshot_id_       ( cflow$dflow_snapshot_id_ ),
    .reset                    ( cflow$reset ),
    .commit_status            ( cflow$commit_status ),
    .register_serialize       ( cflow$register_serialize ),
    .dflow_snapshot_rdy       ( cflow$dflow_snapshot_rdy ),
    .check_kill_kill          ( cflow$check_kill_kill ),
    .dflow_free_snapshot_id_  ( cflow$dflow_free_snapshot_id_ ),
    .dflow_restore_source_id  ( cflow$dflow_restore_source_id ),
    .get_head_seq             ( cflow$get_head_seq ),
    .register_success         ( cflow$register_success ),
    .dflow_rollback_call      ( cflow$dflow_rollback_call ),
    .dflow_snapshot_call      ( cflow$dflow_snapshot_call ),
    .register_spec_idx        ( cflow$register_spec_idx ),
    .check_redirect_target    ( cflow$check_redirect_target ),
    .dflow_free_snapshot_call ( cflow$dflow_free_snapshot_call ),
    .check_redirect_redirect  ( cflow$check_redirect_redirect ),
    .get_head_rdy             ( cflow$get_head_rdy ),
    .register_branch_mask     ( cflow$register_branch_mask ),
    .dflow_restore_call       ( cflow$dflow_restore_call ),
    .register_seq             ( cflow$register_seq )
  );

  // commit temporaries
  logic   [   0:0] commit$cflow_get_head_rdy;
  logic   [ 141:0] commit$in_peek_msg;
  logic   [   0:0] commit$clk;
  logic   [   4:0] commit$kill_notify_msg;
  logic   [   0:0] commit$in_peek_rdy;
  logic   [   3:0] commit$cflow_get_head_seq;
  logic   [   0:0] commit$reset;
  logic   [   1:0] commit$cflow_commit_status;
  logic   [   5:0] commit$dataflow_commit_tag;
  logic   [   0:0] commit$in_take_call;
  logic   [   0:0] commit$dataflow_commit_call;
  logic   [   0:0] commit$cflow_commit_call;

  Commit_0x7d8cae7cdd7a2d86 commit
  (
    .cflow_get_head_rdy   ( commit$cflow_get_head_rdy ),
    .in_peek_msg          ( commit$in_peek_msg ),
    .clk                  ( commit$clk ),
    .kill_notify_msg      ( commit$kill_notify_msg ),
    .in_peek_rdy          ( commit$in_peek_rdy ),
    .cflow_get_head_seq   ( commit$cflow_get_head_seq ),
    .reset                ( commit$reset ),
    .cflow_commit_status  ( commit$cflow_commit_status ),
    .dataflow_commit_tag  ( commit$dataflow_commit_tag ),
    .in_take_call         ( commit$in_take_call ),
    .dataflow_commit_call ( commit$dataflow_commit_call ),
    .cflow_commit_call    ( commit$cflow_commit_call )
  );

  // fetch temporaries
  logic   [  75:0] fetch$mem_recv_msg;
  logic   [   0:0] fetch$clk;
  logic   [   0:0] fetch$mem_recv_rdy;
  logic   [  63:0] fetch$check_redirect_target;
  logic   [   0:0] fetch$reset;
  logic   [   0:0] fetch$take_call;
  logic   [   0:0] fetch$mem_send_rdy;
  logic   [   0:0] fetch$check_redirect_redirect;
  logic   [ 161:0] fetch$peek_msg;
  logic   [ 135:0] fetch$mem_send_msg;
  logic   [   0:0] fetch$peek_rdy;
  logic   [   0:0] fetch$mem_send_call;
  logic   [   0:0] fetch$mem_recv_call;

  Fetch_0x4aa1acfe24534b0 fetch
  (
    .mem_recv_msg            ( fetch$mem_recv_msg ),
    .clk                     ( fetch$clk ),
    .mem_recv_rdy            ( fetch$mem_recv_rdy ),
    .check_redirect_target   ( fetch$check_redirect_target ),
    .reset                   ( fetch$reset ),
    .take_call               ( fetch$take_call ),
    .mem_send_rdy            ( fetch$mem_send_rdy ),
    .check_redirect_redirect ( fetch$check_redirect_redirect ),
    .peek_msg                ( fetch$peek_msg ),
    .mem_send_msg            ( fetch$mem_send_msg ),
    .peek_rdy                ( fetch$peek_rdy ),
    .mem_send_call           ( fetch$mem_send_call ),
    .mem_recv_call           ( fetch$mem_recv_call )
  );

  // signal connections
  assign alu$clk                                   = clk;
  assign alu$in_peek_msg                           = pipe_selector$alu_peek_msg;
  assign alu$in_peek_rdy                           = pipe_selector$alu_peek_rdy;
  assign alu$kill_notify_msg                       = kill_notifier$kill_notify_msg;
  assign alu$reset                                 = reset;
  assign alu$take_call                             = writeback_arbiter$alu_take_call;
  assign branch$clk                                = clk;
  assign branch$in_peek_msg                        = pipe_selector$branch_peek_msg;
  assign branch$in_peek_rdy                        = pipe_selector$branch_peek_rdy;
  assign branch$reset                              = reset;
  assign branch$take_call                          = writeback_arbiter$branch_take_call;
  assign cflow$clk                                 = clk;
  assign cflow$commit_call                         = commit$cflow_commit_call;
  assign cflow$commit_status                       = commit$cflow_commit_status;
  assign cflow$dflow_snapshot_id_                  = dflow$snapshot_id_;
  assign cflow$dflow_snapshot_rdy                  = dflow$snapshot_rdy;
  assign cflow$redirect_call                       = branch$cflow_redirect_call;
  assign cflow$redirect_force                      = branch$cflow_redirect_force;
  assign cflow$redirect_seq                        = branch$cflow_redirect_seq;
  assign cflow$redirect_spec_idx                   = branch$cflow_redirect_spec_idx;
  assign cflow$redirect_target                     = branch$cflow_redirect_target;
  assign cflow$register_call                       = rename$register_call;
  assign cflow$register_pc                         = rename$register_pc;
  assign cflow$register_pc_succ                    = rename$register_pc_succ;
  assign cflow$register_serialize                  = rename$register_serialize;
  assign cflow$register_speculative                = rename$register_speculative;
  assign cflow$reset                               = reset;
  assign commit$cflow_get_head_rdy                 = cflow$get_head_rdy;
  assign commit$cflow_get_head_seq                 = cflow$get_head_seq;
  assign commit$clk                                = clk;
  assign commit$in_peek_msg                        = writeback$peek_msg;
  assign commit$in_peek_rdy                        = writeback$peek_rdy;
  assign commit$kill_notify_msg                    = kill_notifier$kill_notify_msg;
  assign commit$reset                              = reset;
  assign csr$clk                                   = clk;
  assign csr$debug_recv_msg                        = db_recv_msg;
  assign csr$debug_recv_rdy                        = db_recv_rdy;
  assign csr$debug_send_rdy                        = db_send_rdy;
  assign csr$op_call                               = csr_pipe$csr_op_call;
  assign csr$op_csr                                = csr_pipe$csr_op_csr;
  assign csr$op_op                                 = csr_pipe$csr_op_op;
  assign csr$op_rs1_is_x0                          = csr_pipe$csr_op_rs1_is_x0;
  assign csr$op_value                              = csr_pipe$csr_op_value;
  assign csr$reset                                 = reset;
  assign csr_pipe$clk                              = clk;
  assign csr_pipe$csr_op_old                       = csr$op_old;
  assign csr_pipe$csr_op_success                   = csr$op_success;
  assign csr_pipe$in_peek_msg                      = pipe_selector$csr_peek_msg;
  assign csr_pipe$in_peek_rdy                      = pipe_selector$csr_peek_rdy;
  assign csr_pipe$kill_notify_msg                  = kill_notifier$kill_notify_msg;
  assign csr_pipe$reset                            = reset;
  assign csr_pipe$take_call                        = writeback_arbiter$csr_take_call;
  assign db_recv_call                              = csr$debug_recv_call;
  assign db_send_call                              = csr$debug_send_call;
  assign db_send_msg                               = csr$debug_send_msg;
  assign decode$clk                                = clk;
  assign decode$in_peek_msg                        = fetch$peek_msg;
  assign decode$in_peek_rdy                        = fetch$peek_rdy;
  assign decode$kill_notify_msg                    = redirect_notifier$kill_notify_msg;
  assign decode$reset                              = reset;
  assign decode$take_call                          = rename$in_take_call;
  assign dflow$clk                                 = clk;
  assign dflow$commit_call$000                     = commit$dataflow_commit_call;
  assign dflow$commit_tag$000                      = commit$dataflow_commit_tag;
  assign dflow$free_snapshot_call                  = cflow$dflow_free_snapshot_call;
  assign dflow$free_snapshot_id_                   = cflow$dflow_free_snapshot_id_;
  assign dflow$get_dst_areg$000                    = rename$get_dst_areg;
  assign dflow$get_dst_call$000                    = rename$get_dst_call;
  assign dflow$get_src_areg$000                    = rename$get_src_areg$000;
  assign dflow$get_src_areg$001                    = rename$get_src_areg$001;
  assign dflow$is_ready_tag$000                    = issue$is_ready_tag$000;
  assign dflow$is_ready_tag$001                    = issue$is_ready_tag$001;
  assign dflow$read_tag$000                        = dispatch$read_tag$000;
  assign dflow$read_tag$001                        = dispatch$read_tag$001;
  assign dflow$reset                               = reset;
  assign dflow$restore_call                        = cflow$dflow_restore_call;
  assign dflow$restore_source_id                   = cflow$dflow_restore_source_id;
  assign dflow$rollback_call                       = cflow$dflow_rollback_call;
  assign dflow$snapshot_call                       = cflow$dflow_snapshot_call;
  assign dflow$write_call$000                      = writeback$dataflow_write_call;
  assign dflow$write_tag$000                       = writeback$dataflow_write_tag;
  assign dflow$write_value$000                     = writeback$dataflow_write_value;
  assign dispatch$clk                              = clk;
  assign dispatch$in_peek_msg                      = issue$peek_msg;
  assign dispatch$in_peek_rdy                      = issue$peek_rdy;
  assign dispatch$kill_notify_msg                  = kill_notifier$kill_notify_msg;
  assign dispatch$read_value$000                   = dflow$read_value$000;
  assign dispatch$read_value$001                   = dflow$read_value$001;
  assign dispatch$reset                            = reset;
  assign dispatch$take_call                        = pipe_selector$in_take_call;
  assign fetch$check_redirect_redirect             = cflow$check_redirect_redirect;
  assign fetch$check_redirect_target               = cflow$check_redirect_target;
  assign fetch$clk                                 = clk;
  assign fetch$mem_recv_msg                        = mb_recv_0_msg;
  assign fetch$mem_recv_rdy                        = mb_recv_0_rdy;
  assign fetch$mem_send_rdy                        = mb_send_0_rdy;
  assign fetch$reset                               = reset;
  assign fetch$take_call                           = decode$in_take_call;
  assign issue$clk                                 = clk;
  assign issue$get_updated_mask                    = dflow$get_updated_mask;
  assign issue$in_peek_msg                         = rename$peek_msg;
  assign issue$in_peek_rdy                         = rename$peek_rdy;
  assign issue$is_ready_ready$000                  = dflow$is_ready_ready$000;
  assign issue$is_ready_ready$001                  = dflow$is_ready_ready$001;
  assign issue$kill_notify_msg                     = kill_notifier$kill_notify_msg;
  assign issue$reset                               = reset;
  assign issue$take_call                           = dispatch$in_take_call;
  assign kill_notifier$check_kill_kill             = cflow$check_kill_kill;
  assign kill_notifier$clk                         = clk;
  assign kill_notifier$reset                       = reset;
  assign mb_recv_0_call                            = fetch$mem_recv_call;
  assign mb_send_0_call                            = fetch$mem_send_call;
  assign mb_send_0_msg                             = fetch$mem_send_msg;
  assign pipe_selector$alu_take_call               = alu$in_take_call;
  assign pipe_selector$branch_take_call            = branch$in_take_call;
  assign pipe_selector$clk                         = clk;
  assign pipe_selector$csr_take_call               = csr_pipe$in_take_call;
  assign pipe_selector$in_peek_msg                 = dispatch$peek_msg;
  assign pipe_selector$in_peek_rdy                 = dispatch$peek_rdy;
  assign pipe_selector$reset                       = reset;
  assign redirect_notifier$check_redirect_redirect = cflow$check_redirect_redirect;
  assign redirect_notifier$check_redirect_target   = cflow$check_redirect_target;
  assign redirect_notifier$clk                     = clk;
  assign redirect_notifier$reset                   = reset;
  assign rename$clk                                = clk;
  assign rename$get_dst_preg                       = dflow$get_dst_preg$000;
  assign rename$get_dst_rdy                        = dflow$get_dst_rdy$000;
  assign rename$get_src_preg$000                   = dflow$get_src_preg$000;
  assign rename$get_src_preg$001                   = dflow$get_src_preg$001;
  assign rename$in_peek_msg                        = decode$peek_msg;
  assign rename$in_peek_rdy                        = decode$peek_rdy;
  assign rename$kill_notify_msg                    = kill_notifier$kill_notify_msg;
  assign rename$register_branch_mask               = cflow$register_branch_mask;
  assign rename$register_seq                       = cflow$register_seq;
  assign rename$register_spec_idx                  = cflow$register_spec_idx;
  assign rename$register_success                   = cflow$register_success;
  assign rename$reset                              = reset;
  assign rename$take_call                          = issue$in_take_call;
  assign writeback$clk                             = clk;
  assign writeback$in_peek_msg                     = writeback_arbiter$peek_msg;
  assign writeback$in_peek_rdy                     = writeback_arbiter$peek_rdy;
  assign writeback$kill_notify_msg                 = kill_notifier$kill_notify_msg;
  assign writeback$reset                           = reset;
  assign writeback$take_call                       = commit$in_take_call;
  assign writeback_arbiter$alu_peek_msg            = alu$peek_msg;
  assign writeback_arbiter$alu_peek_rdy            = alu$peek_rdy;
  assign writeback_arbiter$branch_peek_msg         = branch$peek_msg;
  assign writeback_arbiter$branch_peek_rdy         = branch$peek_rdy;
  assign writeback_arbiter$clk                     = clk;
  assign writeback_arbiter$csr_peek_msg            = csr_pipe$peek_msg;
  assign writeback_arbiter$csr_peek_rdy            = csr_pipe$peek_rdy;
  assign writeback_arbiter$reset                   = reset;
  assign writeback_arbiter$take_call               = writeback$in_take_call;



endmodule // proc

//-----------------------------------------------------------------------------
// GS11LRenameStage20LRenameDropController_0x6f71125cae5ffc5
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"args": ["process <C> (in_: Bits(190)) -> (accepted: Bits(1), out: Bits(142))"], "kwargs": {}}
// PyMTL: verilator_xinit = zeros
module GS11LRenameStage20LRenameDropController_0x6f71125cae5ffc5
(
  input  logic [   0:0] clk,
  output logic [   4:0] get_dst_areg,
  output logic [   0:0] get_dst_call,
  input  logic [   5:0] get_dst_preg,
  input  logic [   0:0] get_dst_rdy,
  output logic [   4:0] get_src_areg$000,
  output logic [   4:0] get_src_areg$001,
  input  logic [   5:0] get_src_preg$000,
  input  logic [   5:0] get_src_preg$001,
  input  logic [ 189:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 141:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   1:0] register_branch_mask,
  output logic [   0:0] register_call,
  output logic [  63:0] register_pc,
  output logic [  63:0] register_pc_succ,
  input  logic [   3:0] register_seq,
  output logic [   0:0] register_serialize,
  input  logic [   0:0] register_spec_idx,
  output logic [   0:0] register_speculative,
  input  logic [   0:0] register_success,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // pipeline_stage temporaries
  logic   [   0:0] pipeline_stage$check_keep;
  logic   [ 189:0] pipeline_stage$in_peek_msg;
  logic   [   0:0] pipeline_stage$clk;
  logic   [   4:0] pipeline_stage$kill_notify_msg;
  logic   [   0:0] pipeline_stage$in_peek_rdy;
  logic   [   0:0] pipeline_stage$process_accepted;
  logic   [ 141:0] pipeline_stage$check_out;
  logic   [   0:0] pipeline_stage$reset;
  logic   [ 141:0] pipeline_stage$process_out;
  logic   [   0:0] pipeline_stage$take_call;
  logic   [   0:0] pipeline_stage$process_call;
  logic   [ 141:0] pipeline_stage$check_in_;
  logic   [ 141:0] pipeline_stage$peek_msg;
  logic   [   4:0] pipeline_stage$check_msg;
  logic   [   0:0] pipeline_stage$in_take_call;
  logic   [   0:0] pipeline_stage$peek_rdy;
  logic   [ 189:0] pipeline_stage$process_in_;

  PipelineStage_0x66dba493805010c7 pipeline_stage
  (
    .check_keep       ( pipeline_stage$check_keep ),
    .in_peek_msg      ( pipeline_stage$in_peek_msg ),
    .clk              ( pipeline_stage$clk ),
    .kill_notify_msg  ( pipeline_stage$kill_notify_msg ),
    .in_peek_rdy      ( pipeline_stage$in_peek_rdy ),
    .process_accepted ( pipeline_stage$process_accepted ),
    .check_out        ( pipeline_stage$check_out ),
    .reset            ( pipeline_stage$reset ),
    .process_out      ( pipeline_stage$process_out ),
    .take_call        ( pipeline_stage$take_call ),
    .process_call     ( pipeline_stage$process_call ),
    .check_in_        ( pipeline_stage$check_in_ ),
    .peek_msg         ( pipeline_stage$peek_msg ),
    .check_msg        ( pipeline_stage$check_msg ),
    .in_take_call     ( pipeline_stage$in_take_call ),
    .peek_rdy         ( pipeline_stage$peek_rdy ),
    .process_in_      ( pipeline_stage$process_in_ )
  );

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [ 141:0] drop_controller$check_in_;
  logic   [   4:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [ 141:0] drop_controller$check_out;

  PipelineKillDropController_0x6535c882219b5c15 drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // stage temporaries
  logic   [   5:0] stage$get_dst_preg;
  logic   [   1:0] stage$register_branch_mask;
  logic   [   0:0] stage$process_call;
  logic   [   0:0] stage$clk;
  logic   [   5:0] stage$get_src_preg$000;
  logic   [   5:0] stage$get_src_preg$001;
  logic   [   0:0] stage$get_dst_rdy;
  logic   [   0:0] stage$register_spec_idx;
  logic   [   0:0] stage$reset;
  logic   [   0:0] stage$register_success;
  logic   [ 189:0] stage$process_in_;
  logic   [   3:0] stage$register_seq;
  logic   [   4:0] stage$get_src_areg$000;
  logic   [   4:0] stage$get_src_areg$001;
  logic   [   4:0] stage$get_dst_areg;
  logic   [   0:0] stage$process_accepted;
  logic   [  63:0] stage$register_pc;
  logic   [   0:0] stage$register_speculative;
  logic   [   0:0] stage$get_dst_call;
  logic   [   0:0] stage$register_call;
  logic   [   0:0] stage$register_serialize;
  logic   [ 141:0] stage$process_out;
  logic   [  63:0] stage$register_pc_succ;

  RenameStage_0x6ed532e713c6d3 stage
  (
    .get_dst_preg         ( stage$get_dst_preg ),
    .register_branch_mask ( stage$register_branch_mask ),
    .process_call         ( stage$process_call ),
    .clk                  ( stage$clk ),
    .get_src_preg$000     ( stage$get_src_preg$000 ),
    .get_src_preg$001     ( stage$get_src_preg$001 ),
    .get_dst_rdy          ( stage$get_dst_rdy ),
    .register_spec_idx    ( stage$register_spec_idx ),
    .reset                ( stage$reset ),
    .register_success     ( stage$register_success ),
    .process_in_          ( stage$process_in_ ),
    .register_seq         ( stage$register_seq ),
    .get_src_areg$000     ( stage$get_src_areg$000 ),
    .get_src_areg$001     ( stage$get_src_areg$001 ),
    .get_dst_areg         ( stage$get_dst_areg ),
    .process_accepted     ( stage$process_accepted ),
    .register_pc          ( stage$register_pc ),
    .register_speculative ( stage$register_speculative ),
    .get_dst_call         ( stage$get_dst_call ),
    .register_call        ( stage$register_call ),
    .register_serialize   ( stage$register_serialize ),
    .process_out          ( stage$process_out ),
    .register_pc_succ     ( stage$register_pc_succ )
  );

  // signal connections
  assign drop_controller$check_in_       = pipeline_stage$check_in_;
  assign drop_controller$check_msg       = pipeline_stage$check_msg;
  assign drop_controller$clk             = clk;
  assign drop_controller$reset           = reset;
  assign get_dst_areg                    = stage$get_dst_areg;
  assign get_dst_call                    = stage$get_dst_call;
  assign get_src_areg$000                = stage$get_src_areg$000;
  assign get_src_areg$001                = stage$get_src_areg$001;
  assign in_take_call                    = pipeline_stage$in_take_call;
  assign peek_msg                        = pipeline_stage$peek_msg;
  assign peek_rdy                        = pipeline_stage$peek_rdy;
  assign pipeline_stage$check_keep       = drop_controller$check_keep;
  assign pipeline_stage$check_out        = drop_controller$check_out;
  assign pipeline_stage$clk              = clk;
  assign pipeline_stage$in_peek_msg      = in_peek_msg;
  assign pipeline_stage$in_peek_rdy      = in_peek_rdy;
  assign pipeline_stage$kill_notify_msg  = kill_notify_msg;
  assign pipeline_stage$process_accepted = stage$process_accepted;
  assign pipeline_stage$process_out      = stage$process_out;
  assign pipeline_stage$reset            = reset;
  assign pipeline_stage$take_call        = take_call;
  assign register_call                   = stage$register_call;
  assign register_pc                     = stage$register_pc;
  assign register_pc_succ                = stage$register_pc_succ;
  assign register_serialize              = stage$register_serialize;
  assign register_speculative            = stage$register_speculative;
  assign stage$clk                       = clk;
  assign stage$get_dst_preg              = get_dst_preg;
  assign stage$get_dst_rdy               = get_dst_rdy;
  assign stage$get_src_preg$000          = get_src_preg$000;
  assign stage$get_src_preg$001          = get_src_preg$001;
  assign stage$process_call              = pipeline_stage$process_call;
  assign stage$process_in_               = pipeline_stage$process_in_;
  assign stage$register_branch_mask      = register_branch_mask;
  assign stage$register_seq              = register_seq;
  assign stage$register_spec_idx         = register_spec_idx;
  assign stage$register_success          = register_success;
  assign stage$reset                     = reset;



endmodule // GS11LRenameStage20LRenameDropController_0x6f71125cae5ffc5

//-----------------------------------------------------------------------------
// PipelineStage_0x66dba493805010c7
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"In": 190, "Intermediate": null, "interface": "kill_notify (msg: Bits(5)) -> (); peek <R> () -> (msg: Bits(142)); take <C> () -> ()"}
// PyMTL: verilator_xinit = zeros
module PipelineStage_0x66dba493805010c7
(
  output logic [ 141:0] check_in_,
  input  logic [   0:0] check_keep,
  output logic [   4:0] check_msg,
  input  logic [ 141:0] check_out,
  input  logic [   0:0] clk,
  input  logic [ 189:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 141:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] process_accepted,
  output logic [   0:0] process_call,
  output logic [ 189:0] process_in_,
  input  logic [ 141:0] process_out,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // logic declarations
  logic   [   0:0] output_clear;
  logic   [   0:0] input_available;


  // register declarations
  logic    [   0:0] advance;
  logic    [   0:0] taking;

  // vvm temporaries
  logic   [   0:0] vvm$check_keep;
  logic   [   0:0] vvm$clk;
  logic   [   4:0] vvm$kill_notify_msg;
  logic   [ 141:0] vvm$add_msg;
  logic   [ 141:0] vvm$check_out;
  logic   [   0:0] vvm$reset;
  logic   [   0:0] vvm$add_call;
  logic   [   0:0] vvm$take_call;
  logic   [ 141:0] vvm$check_in_;
  logic   [ 141:0] vvm$peek_msg;
  logic   [   0:0] vvm$add_rdy;
  logic   [   4:0] vvm$check_msg;
  logic   [   0:0] vvm$peek_rdy;

  ValidValueManager_0xed9504a4389a8c9 vvm
  (
    .check_keep      ( vvm$check_keep ),
    .clk             ( vvm$clk ),
    .kill_notify_msg ( vvm$kill_notify_msg ),
    .add_msg         ( vvm$add_msg ),
    .check_out       ( vvm$check_out ),
    .reset           ( vvm$reset ),
    .add_call        ( vvm$add_call ),
    .take_call       ( vvm$take_call ),
    .check_in_       ( vvm$check_in_ ),
    .peek_msg        ( vvm$peek_msg ),
    .add_rdy         ( vvm$add_rdy ),
    .check_msg       ( vvm$check_msg ),
    .peek_rdy        ( vvm$peek_rdy )
  );

  // signal connections
  assign check_in_           = vvm$check_in_;
  assign check_msg           = vvm$check_msg;
  assign in_take_call        = taking;
  assign input_available     = in_peek_rdy;
  assign output_clear        = vvm$add_rdy;
  assign peek_msg            = vvm$peek_msg;
  assign peek_rdy            = vvm$peek_rdy;
  assign process_call        = advance;
  assign process_in_         = in_peek_msg;
  assign vvm$add_call        = taking;
  assign vvm$add_msg         = process_out;
  assign vvm$check_keep      = check_keep;
  assign vvm$check_out       = check_out;
  assign vvm$clk             = clk;
  assign vvm$kill_notify_msg = kill_notify_msg;
  assign vvm$reset           = reset;
  assign vvm$take_call       = take_call;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_taking():
  //       s.taking.v = s.advance & s.process_accepted

  // logic for handle_taking()
  always @ (*) begin
    taking = (advance&process_accepted);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_advance():
  //       s.advance.v = s.output_clear and s.input_available

  // logic for handle_advance()
  always @ (*) begin
    advance = (output_clear&&input_available);
  end


endmodule // PipelineStage_0x66dba493805010c7

//-----------------------------------------------------------------------------
// ValidValueManager_0xed9504a4389a8c9
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"interface": "kill_notify (msg: Bits(5)) -> (); peek <R> () -> (msg: Bits(142)); take <C> () -> (); add <CR> (msg: Bits(142)) -> ()"}
// PyMTL: verilator_xinit = zeros
module ValidValueManager_0xed9504a4389a8c9
(
  input  logic [   0:0] add_call,
  input  logic [ 141:0] add_msg,
  output logic [   0:0] add_rdy,
  output logic [ 141:0] check_in_,
  input  logic [   0:0] check_keep,
  output logic [   4:0] check_msg,
  input  logic [ 141:0] check_out,
  input  logic [   0:0] clk,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 141:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // register declarations
  logic    [   0:0] output_clear;
  logic    [   0:0] output_rdy;
  logic    [   0:0] val_reg$write_data;

  // val_reg temporaries
  logic   [   0:0] val_reg$clk;
  logic   [   0:0] val_reg$reset;
  logic   [   0:0] val_reg$read_data;

  Register_0x360ff20b8ea9d7d7 val_reg
  (
    .clk        ( val_reg$clk ),
    .write_data ( val_reg$write_data ),
    .reset      ( val_reg$reset ),
    .read_data  ( val_reg$read_data )
  );

  // out_reg temporaries
  logic   [   0:0] out_reg$clk;
  logic   [   0:0] out_reg$write_call;
  logic   [ 141:0] out_reg$write_data;
  logic   [   0:0] out_reg$reset;
  logic   [ 141:0] out_reg$read_data;

  Register_0x24d6bb878320116e out_reg
  (
    .clk        ( out_reg$clk ),
    .write_call ( out_reg$write_call ),
    .write_data ( out_reg$write_data ),
    .reset      ( out_reg$reset ),
    .read_data  ( out_reg$read_data )
  );

  // signal connections
  assign add_rdy            = output_clear;
  assign check_in_          = out_reg$read_data;
  assign check_msg          = kill_notify_msg;
  assign out_reg$clk        = clk;
  assign out_reg$reset      = reset;
  assign out_reg$write_call = add_call;
  assign out_reg$write_data = add_msg;
  assign peek_msg           = check_out;
  assign peek_rdy           = output_rdy;
  assign val_reg$clk        = clk;
  assign val_reg$reset      = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_rdy():
  //       if s.val_reg.read_data:
  //         s.output_rdy.v = s.check_keep
  //       else:
  //         s.output_rdy.v = 0

  // logic for handle_rdy()
  always @ (*) begin
    if (val_reg$read_data) begin
      output_rdy = check_keep;
    end
    else begin
      output_rdy = 0;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_clear():
  //       s.output_clear.v = not s.output_rdy or s.take_call

  // logic for handle_clear()
  always @ (*) begin
    output_clear = (!output_rdy||take_call);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_val_reg_in():
  //       if s.add_call:
  //         s.val_reg.write_data.v = 1
  //       else:
  //         s.val_reg.write_data.v = not s.output_clear

  // logic for handle_val_reg_in()
  always @ (*) begin
    if (add_call) begin
      val_reg$write_data = 1;
    end
    else begin
      val_reg$write_data = !output_clear;
    end
  end


endmodule // ValidValueManager_0xed9504a4389a8c9

//-----------------------------------------------------------------------------
// Register_0x360ff20b8ea9d7d7
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(1)); write (data: Bits(1)) -> ()", "reset_value": 0}
// PyMTL: verilator_xinit = zeros
module Register_0x360ff20b8ea9d7d7
(
  input  logic [   0:0] clk,
  output logic [   0:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [   0:0] reg_value;

  // localparam declarations
  localparam reset_value = 0;

  // signal connections
  assign read_data = reg_value;
  assign update    = 1'd1;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.reset:
  //           s.reg_value.n = reset_value
  //         elif s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      reg_value <= reset_value;
    end
    else begin
      if (update) begin
        reg_value <= write_data;
      end
      else begin
      end
    end
  end


endmodule // Register_0x360ff20b8ea9d7d7

//-----------------------------------------------------------------------------
// Register_0x24d6bb878320116e
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(142)); write <C> (data: Bits(142)) -> ()", "reset_value": null}
// PyMTL: verilator_xinit = zeros
module Register_0x24d6bb878320116e
(
  input  logic [   0:0] clk,
  output logic [ 141:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [ 141:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [ 141:0] reg_value;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (update) begin
      reg_value <= write_data;
    end
    else begin
    end
  end


endmodule // Register_0x24d6bb878320116e

//-----------------------------------------------------------------------------
// PipelineKillDropController_0x6535c882219b5c15
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.kill_unit {"interface": "check (msg: Bits(5), in_: Bits(142)) -> (out: Bits(142), keep: Bits(1))"}
// PyMTL: verilator_xinit = zeros
module PipelineKillDropController_0x6535c882219b5c15
(
  input  logic [ 141:0] check_in_,
  output logic [   0:0] check_keep,
  input  logic [   4:0] check_msg,
  output logic  [ 141:0] check_out,
  input  logic [   0:0] clk,
  input  logic [   0:0] reset
);

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [   1:0] drop_controller$check_in_;
  logic   [   4:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [   1:0] drop_controller$check_out;

  KillDropController_0xccf15b584e8c1d drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // signal connections
  assign check_keep                = drop_controller$check_keep;
  assign drop_controller$check_in_ = check_in_[73:72];
  assign drop_controller$check_msg = check_msg;
  assign drop_controller$clk       = clk;
  assign drop_controller$reset     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_out():
  //       # Set the out equal to the input and then override the branch mask
  //       s.check_out.v = s.check_in_
  //       s.check_out.hdr_branch_mask.v = s.drop_controller.check_out

  // logic for handle_out()
  always @ (*) begin
    check_out = check_in_;
    check_out[(74)-1:72] = drop_controller$check_out;
  end


endmodule // PipelineKillDropController_0x6535c882219b5c15

//-----------------------------------------------------------------------------
// KillDropController_0xccf15b584e8c1d
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.kill_unit {"interface": "check (msg: Bits(5), in_: Bits(2)) -> (out: Bits(2), keep: Bits(1))"}
// PyMTL: verilator_xinit = zeros
module KillDropController_0xccf15b584e8c1d
(
  input  logic [   1:0] check_in_,
  output logic  [   0:0] check_keep,
  input  logic [   4:0] check_msg,
  output logic  [   1:0] check_out,
  input  logic [   0:0] clk,
  input  logic [   0:0] reset
);

  // register declarations
  logic    [   1:0] kill_match;



  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_check():
  //       s.kill_match.v = s.check_in_ & s.check_msg.kill_mask
  //       s.check_keep.v = not (reduce_or(s.kill_match) or s.check_msg.force)
  //       s.check_out.v = s.check_in_ & (~s.check_msg.clear_mask)

  // logic for handle_check()
  always @ (*) begin
    kill_match = (check_in_&check_msg[(3)-1:1]);
    check_keep = !((|kill_match)||check_msg[(1)-1:0]);
    check_out = (check_in_&~check_msg[(5)-1:3]);
  end


endmodule // KillDropController_0xccf15b584e8c1d

//-----------------------------------------------------------------------------
// RenameStage_0x6ed532e713c6d3
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.backend.rename {"rename_interface": "process <C> (in_: Bits(190)) -> (accepted: Bits(1), out: Bits(142))"}
// PyMTL: verilator_xinit = zeros
module RenameStage_0x6ed532e713c6d3
(
  input  logic [   0:0] clk,
  output logic [   4:0] get_dst_areg,
  output logic  [   0:0] get_dst_call,
  input  logic [   5:0] get_dst_preg,
  input  logic [   0:0] get_dst_rdy,
  output logic [   4:0] get_src_areg$000,
  output logic [   4:0] get_src_areg$001,
  input  logic [   5:0] get_src_preg$000,
  input  logic [   5:0] get_src_preg$001,
  output logic [   0:0] process_accepted,
  input  logic [   0:0] process_call,
  input  logic [ 189:0] process_in_,
  output logic [ 141:0] process_out,
  input  logic [   1:0] register_branch_mask,
  output logic [   0:0] register_call,
  output logic [  63:0] register_pc,
  output logic [  63:0] register_pc_succ,
  input  logic [   3:0] register_seq,
  output logic [   0:0] register_serialize,
  input  logic [   0:0] register_spec_idx,
  output logic [   0:0] register_speculative,
  input  logic [   0:0] register_success,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [ 189:0] decoded_;
  logic   [   0:0] accepted_;


  // register declarations
  logic    [ 141:0] out_;

  // localparam declarations
  localparam PIPELINE_MSG_STATUS_VALID = 2'd0;

  // signal connections
  assign accepted_            = register_success;
  assign decoded_             = process_in_;
  assign get_dst_areg         = decoded_[149:145];
  assign get_src_areg$000     = decoded_[137:133];
  assign get_src_areg$001     = decoded_[143:139];
  assign process_accepted     = accepted_;
  assign process_out          = out_;
  assign register_call        = process_call;
  assign register_pc          = decoded_[65:2];
  assign register_pc_succ     = decoded_[131:68];
  assign register_serialize   = decoded_[66:66];
  assign register_speculative = decoded_[67:67];

  // array declarations
  logic   [   5:0] get_src_preg[0:1];
  assign get_src_preg[  0] = get_src_preg$000;
  assign get_src_preg[  1] = get_src_preg$001;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_calls():
  //       s.get_dst_call.v = s.accepted_ and s.decoded_.rd_val and (
  //           s.decoded_.hdr_status == PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID)

  // logic for handle_calls()
  always @ (*) begin
    get_dst_call = (accepted_&&decoded_[(145)-1:144]&&(decoded_[(2)-1:0] == PIPELINE_MSG_STATUS_VALID));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_out():
  //       s.out_.v = 0  # No inferred latches
  //       s.out_.hdr_frontend_hdr.v = s.decoded_.hdr
  //       s.out_.hdr_seq.v = s.register_seq
  //       s.out_.hdr_branch_mask.v = s.register_branch_mask
  //       s.out_.hdr_spec_val.v = s.decoded_.speculative
  //       s.out_.hdr_spec.v = s.register_spec_idx
  //       s.out_.hdr_branch_mask.v = s.register_branch_mask
  //       # We need to propogate exception info
  //       if s.decoded_.hdr_status == PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID:
  //         s.out_.rs1_val.v = s.decoded_.rs1_val
  //         s.out_.rs2_val.v = s.decoded_.rs2_val
  //         s.out_.rd_val.v = s.decoded_.rd_val
  //         # Copy over the aregs
  //         s.out_.rs1.v = s.get_src_preg[0]
  //         s.out_.rs2.v = s.get_src_preg[1]
  //         s.out_.rd.v = s.get_dst_preg
  //         # Copy the execution stuff
  //         s.out_.execution_data.v = s.decoded_.execution_data
  //       else:
  //         s.out_.exception_info.v = s.decoded_.exception_info

  // logic for handle_out()
  always @ (*) begin
    out_ = 0;
    out_[(66)-1:0] = decoded_[(66)-1:0];
    out_[(70)-1:66] = register_seq;
    out_[(74)-1:72] = register_branch_mask;
    out_[(71)-1:70] = decoded_[(68)-1:67];
    out_[(72)-1:71] = register_spec_idx;
    out_[(74)-1:72] = register_branch_mask;
    if ((decoded_[(2)-1:0] == PIPELINE_MSG_STATUS_VALID)) begin
      out_[(75)-1:74] = decoded_[(133)-1:132];
      out_[(82)-1:81] = decoded_[(139)-1:138];
      out_[(89)-1:88] = decoded_[(145)-1:144];
      out_[(81)-1:75] = get_src_preg[0];
      out_[(88)-1:82] = get_src_preg[1];
      out_[(95)-1:89] = get_dst_preg;
      out_[(135)-1:95] = decoded_[(190)-1:150];
    end
    else begin
      out_[(142)-1:74] = decoded_[(134)-1:66];
    end
  end


endmodule // RenameStage_0x6ed532e713c6d3

//-----------------------------------------------------------------------------
// GS13LDispatchStage22LDispatchDropController_0x78e60f5988db2eb3
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"args": ["process <C> (in_: Bits(142)) -> (accepted: Bits(1), out: Bits(251))"], "kwargs": {}}
// PyMTL: verilator_xinit = zeros
module GS13LDispatchStage22LDispatchDropController_0x78e60f5988db2eb3
(
  input  logic [   0:0] clk,
  input  logic [ 141:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 250:0] peek_msg,
  output logic [   0:0] peek_rdy,
  output logic [   5:0] read_tag$000,
  output logic [   5:0] read_tag$001,
  input  logic [  63:0] read_value$000,
  input  logic [  63:0] read_value$001,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // pipeline_stage temporaries
  logic   [   0:0] pipeline_stage$check_keep;
  logic   [ 141:0] pipeline_stage$in_peek_msg;
  logic   [   0:0] pipeline_stage$clk;
  logic   [   4:0] pipeline_stage$kill_notify_msg;
  logic   [   0:0] pipeline_stage$in_peek_rdy;
  logic   [   0:0] pipeline_stage$process_accepted;
  logic   [ 250:0] pipeline_stage$check_out;
  logic   [   0:0] pipeline_stage$reset;
  logic   [ 250:0] pipeline_stage$process_out;
  logic   [   0:0] pipeline_stage$take_call;
  logic   [   0:0] pipeline_stage$process_call;
  logic   [ 250:0] pipeline_stage$check_in_;
  logic   [ 250:0] pipeline_stage$peek_msg;
  logic   [   4:0] pipeline_stage$check_msg;
  logic   [   0:0] pipeline_stage$in_take_call;
  logic   [   0:0] pipeline_stage$peek_rdy;
  logic   [ 141:0] pipeline_stage$process_in_;

  PipelineStage_0x1289115dcfdf81a7 pipeline_stage
  (
    .check_keep       ( pipeline_stage$check_keep ),
    .in_peek_msg      ( pipeline_stage$in_peek_msg ),
    .clk              ( pipeline_stage$clk ),
    .kill_notify_msg  ( pipeline_stage$kill_notify_msg ),
    .in_peek_rdy      ( pipeline_stage$in_peek_rdy ),
    .process_accepted ( pipeline_stage$process_accepted ),
    .check_out        ( pipeline_stage$check_out ),
    .reset            ( pipeline_stage$reset ),
    .process_out      ( pipeline_stage$process_out ),
    .take_call        ( pipeline_stage$take_call ),
    .process_call     ( pipeline_stage$process_call ),
    .check_in_        ( pipeline_stage$check_in_ ),
    .peek_msg         ( pipeline_stage$peek_msg ),
    .check_msg        ( pipeline_stage$check_msg ),
    .in_take_call     ( pipeline_stage$in_take_call ),
    .peek_rdy         ( pipeline_stage$peek_rdy ),
    .process_in_      ( pipeline_stage$process_in_ )
  );

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [ 250:0] drop_controller$check_in_;
  logic   [   4:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [ 250:0] drop_controller$check_out;

  PipelineKillDropController_0x7f2faca09c5dd2f7 drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // stage temporaries
  logic   [   0:0] stage$process_call;
  logic   [   0:0] stage$clk;
  logic   [  63:0] stage$read_value$000;
  logic   [  63:0] stage$read_value$001;
  logic   [   0:0] stage$reset;
  logic   [ 141:0] stage$process_in_;
  logic   [   0:0] stage$process_accepted;
  logic   [   5:0] stage$read_tag$000;
  logic   [   5:0] stage$read_tag$001;
  logic   [ 250:0] stage$process_out;

  DispatchStage_0x3d3671bf74513fd9 stage
  (
    .process_call     ( stage$process_call ),
    .clk              ( stage$clk ),
    .read_value$000   ( stage$read_value$000 ),
    .read_value$001   ( stage$read_value$001 ),
    .reset            ( stage$reset ),
    .process_in_      ( stage$process_in_ ),
    .process_accepted ( stage$process_accepted ),
    .read_tag$000     ( stage$read_tag$000 ),
    .read_tag$001     ( stage$read_tag$001 ),
    .process_out      ( stage$process_out )
  );

  // signal connections
  assign drop_controller$check_in_       = pipeline_stage$check_in_;
  assign drop_controller$check_msg       = pipeline_stage$check_msg;
  assign drop_controller$clk             = clk;
  assign drop_controller$reset           = reset;
  assign in_take_call                    = pipeline_stage$in_take_call;
  assign peek_msg                        = pipeline_stage$peek_msg;
  assign peek_rdy                        = pipeline_stage$peek_rdy;
  assign pipeline_stage$check_keep       = drop_controller$check_keep;
  assign pipeline_stage$check_out        = drop_controller$check_out;
  assign pipeline_stage$clk              = clk;
  assign pipeline_stage$in_peek_msg      = in_peek_msg;
  assign pipeline_stage$in_peek_rdy      = in_peek_rdy;
  assign pipeline_stage$kill_notify_msg  = kill_notify_msg;
  assign pipeline_stage$process_accepted = stage$process_accepted;
  assign pipeline_stage$process_out      = stage$process_out;
  assign pipeline_stage$reset            = reset;
  assign pipeline_stage$take_call        = take_call;
  assign read_tag$000                    = stage$read_tag$000;
  assign read_tag$001                    = stage$read_tag$001;
  assign stage$clk                       = clk;
  assign stage$process_call              = pipeline_stage$process_call;
  assign stage$process_in_               = pipeline_stage$process_in_;
  assign stage$read_value$000            = read_value$000;
  assign stage$read_value$001            = read_value$001;
  assign stage$reset                     = reset;



endmodule // GS13LDispatchStage22LDispatchDropController_0x78e60f5988db2eb3

//-----------------------------------------------------------------------------
// PipelineStage_0x1289115dcfdf81a7
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"In": 142, "Intermediate": null, "interface": "kill_notify (msg: Bits(5)) -> (); peek <R> () -> (msg: Bits(251)); take <C> () -> ()"}
// PyMTL: verilator_xinit = zeros
module PipelineStage_0x1289115dcfdf81a7
(
  output logic [ 250:0] check_in_,
  input  logic [   0:0] check_keep,
  output logic [   4:0] check_msg,
  input  logic [ 250:0] check_out,
  input  logic [   0:0] clk,
  input  logic [ 141:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 250:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] process_accepted,
  output logic [   0:0] process_call,
  output logic [ 141:0] process_in_,
  input  logic [ 250:0] process_out,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // logic declarations
  logic   [   0:0] output_clear;
  logic   [   0:0] input_available;


  // register declarations
  logic    [   0:0] advance;
  logic    [   0:0] taking;

  // vvm temporaries
  logic   [   0:0] vvm$check_keep;
  logic   [   0:0] vvm$clk;
  logic   [   4:0] vvm$kill_notify_msg;
  logic   [ 250:0] vvm$add_msg;
  logic   [ 250:0] vvm$check_out;
  logic   [   0:0] vvm$reset;
  logic   [   0:0] vvm$add_call;
  logic   [   0:0] vvm$take_call;
  logic   [ 250:0] vvm$check_in_;
  logic   [ 250:0] vvm$peek_msg;
  logic   [   0:0] vvm$add_rdy;
  logic   [   4:0] vvm$check_msg;
  logic   [   0:0] vvm$peek_rdy;

  ValidValueManager_0x369c9400f0e2a885 vvm
  (
    .check_keep      ( vvm$check_keep ),
    .clk             ( vvm$clk ),
    .kill_notify_msg ( vvm$kill_notify_msg ),
    .add_msg         ( vvm$add_msg ),
    .check_out       ( vvm$check_out ),
    .reset           ( vvm$reset ),
    .add_call        ( vvm$add_call ),
    .take_call       ( vvm$take_call ),
    .check_in_       ( vvm$check_in_ ),
    .peek_msg        ( vvm$peek_msg ),
    .add_rdy         ( vvm$add_rdy ),
    .check_msg       ( vvm$check_msg ),
    .peek_rdy        ( vvm$peek_rdy )
  );

  // signal connections
  assign check_in_           = vvm$check_in_;
  assign check_msg           = vvm$check_msg;
  assign in_take_call        = taking;
  assign input_available     = in_peek_rdy;
  assign output_clear        = vvm$add_rdy;
  assign peek_msg            = vvm$peek_msg;
  assign peek_rdy            = vvm$peek_rdy;
  assign process_call        = advance;
  assign process_in_         = in_peek_msg;
  assign vvm$add_call        = taking;
  assign vvm$add_msg         = process_out;
  assign vvm$check_keep      = check_keep;
  assign vvm$check_out       = check_out;
  assign vvm$clk             = clk;
  assign vvm$kill_notify_msg = kill_notify_msg;
  assign vvm$reset           = reset;
  assign vvm$take_call       = take_call;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_taking():
  //       s.taking.v = s.advance & s.process_accepted

  // logic for handle_taking()
  always @ (*) begin
    taking = (advance&process_accepted);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_advance():
  //       s.advance.v = s.output_clear and s.input_available

  // logic for handle_advance()
  always @ (*) begin
    advance = (output_clear&&input_available);
  end


endmodule // PipelineStage_0x1289115dcfdf81a7

//-----------------------------------------------------------------------------
// ValidValueManager_0x369c9400f0e2a885
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"interface": "kill_notify (msg: Bits(5)) -> (); peek <R> () -> (msg: Bits(251)); take <C> () -> (); add <CR> (msg: Bits(251)) -> ()"}
// PyMTL: verilator_xinit = zeros
module ValidValueManager_0x369c9400f0e2a885
(
  input  logic [   0:0] add_call,
  input  logic [ 250:0] add_msg,
  output logic [   0:0] add_rdy,
  output logic [ 250:0] check_in_,
  input  logic [   0:0] check_keep,
  output logic [   4:0] check_msg,
  input  logic [ 250:0] check_out,
  input  logic [   0:0] clk,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 250:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // register declarations
  logic    [   0:0] output_clear;
  logic    [   0:0] output_rdy;
  logic    [   0:0] val_reg$write_data;

  // val_reg temporaries
  logic   [   0:0] val_reg$clk;
  logic   [   0:0] val_reg$reset;
  logic   [   0:0] val_reg$read_data;

  Register_0x360ff20b8ea9d7d7 val_reg
  (
    .clk        ( val_reg$clk ),
    .write_data ( val_reg$write_data ),
    .reset      ( val_reg$reset ),
    .read_data  ( val_reg$read_data )
  );

  // out_reg temporaries
  logic   [   0:0] out_reg$clk;
  logic   [   0:0] out_reg$write_call;
  logic   [ 250:0] out_reg$write_data;
  logic   [   0:0] out_reg$reset;
  logic   [ 250:0] out_reg$read_data;

  Register_0x2b6e6e2a5b9fe130 out_reg
  (
    .clk        ( out_reg$clk ),
    .write_call ( out_reg$write_call ),
    .write_data ( out_reg$write_data ),
    .reset      ( out_reg$reset ),
    .read_data  ( out_reg$read_data )
  );

  // signal connections
  assign add_rdy            = output_clear;
  assign check_in_          = out_reg$read_data;
  assign check_msg          = kill_notify_msg;
  assign out_reg$clk        = clk;
  assign out_reg$reset      = reset;
  assign out_reg$write_call = add_call;
  assign out_reg$write_data = add_msg;
  assign peek_msg           = check_out;
  assign peek_rdy           = output_rdy;
  assign val_reg$clk        = clk;
  assign val_reg$reset      = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_rdy():
  //       if s.val_reg.read_data:
  //         s.output_rdy.v = s.check_keep
  //       else:
  //         s.output_rdy.v = 0

  // logic for handle_rdy()
  always @ (*) begin
    if (val_reg$read_data) begin
      output_rdy = check_keep;
    end
    else begin
      output_rdy = 0;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_clear():
  //       s.output_clear.v = not s.output_rdy or s.take_call

  // logic for handle_clear()
  always @ (*) begin
    output_clear = (!output_rdy||take_call);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_val_reg_in():
  //       if s.add_call:
  //         s.val_reg.write_data.v = 1
  //       else:
  //         s.val_reg.write_data.v = not s.output_clear

  // logic for handle_val_reg_in()
  always @ (*) begin
    if (add_call) begin
      val_reg$write_data = 1;
    end
    else begin
      val_reg$write_data = !output_clear;
    end
  end


endmodule // ValidValueManager_0x369c9400f0e2a885

//-----------------------------------------------------------------------------
// Register_0x2b6e6e2a5b9fe130
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(251)); write <C> (data: Bits(251)) -> ()", "reset_value": null}
// PyMTL: verilator_xinit = zeros
module Register_0x2b6e6e2a5b9fe130
(
  input  logic [   0:0] clk,
  output logic [ 250:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [ 250:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [ 250:0] reg_value;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (update) begin
      reg_value <= write_data;
    end
    else begin
    end
  end


endmodule // Register_0x2b6e6e2a5b9fe130

//-----------------------------------------------------------------------------
// PipelineKillDropController_0x7f2faca09c5dd2f7
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.kill_unit {"interface": "check (msg: Bits(5), in_: Bits(251)) -> (out: Bits(251), keep: Bits(1))"}
// PyMTL: verilator_xinit = zeros
module PipelineKillDropController_0x7f2faca09c5dd2f7
(
  input  logic [ 250:0] check_in_,
  output logic [   0:0] check_keep,
  input  logic [   4:0] check_msg,
  output logic  [ 250:0] check_out,
  input  logic [   0:0] clk,
  input  logic [   0:0] reset
);

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [   1:0] drop_controller$check_in_;
  logic   [   4:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [   1:0] drop_controller$check_out;

  KillDropController_0xccf15b584e8c1d drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // signal connections
  assign check_keep                = drop_controller$check_keep;
  assign drop_controller$check_in_ = check_in_[73:72];
  assign drop_controller$check_msg = check_msg;
  assign drop_controller$clk       = clk;
  assign drop_controller$reset     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_out():
  //       # Set the out equal to the input and then override the branch mask
  //       s.check_out.v = s.check_in_
  //       s.check_out.hdr_branch_mask.v = s.drop_controller.check_out

  // logic for handle_out()
  always @ (*) begin
    check_out = check_in_;
    check_out[(74)-1:72] = drop_controller$check_out;
  end


endmodule // PipelineKillDropController_0x7f2faca09c5dd2f7

//-----------------------------------------------------------------------------
// DispatchStage_0x3d3671bf74513fd9
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.backend.dispatch {"dispatch_interface": "process <C> (in_: Bits(142)) -> (accepted: Bits(1), out: Bits(251))"}
// PyMTL: verilator_xinit = zeros
module DispatchStage_0x3d3671bf74513fd9
(
  input  logic [   0:0] clk,
  output logic [   0:0] process_accepted,
  input  logic [   0:0] process_call,
  input  logic [ 141:0] process_in_,
  output logic [ 250:0] process_out,
  output logic [   5:0] read_tag$000,
  output logic [   5:0] read_tag$001,
  input  logic [  63:0] read_value$000,
  input  logic [  63:0] read_value$001,
  input  logic [   0:0] reset
);

  // register declarations
  logic    [ 250:0] dispatched_;

  // localparam declarations
  localparam PIPELINE_MSG_STATUS_VALID = 2'd0;

  // signal connections
  assign process_accepted = 1'd1;
  assign process_out      = dispatched_;
  assign read_tag$000     = process_in_[80:75];
  assign read_tag$001     = process_in_[87:82];

  // array declarations
  logic   [  63:0] read_value[0:1];
  assign read_value[  0] = read_value$000;
  assign read_value[  1] = read_value$001;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_output():
  //       s.dispatched_.v = 0
  //       s.dispatched_.hdr.v = s.process_in_.hdr
  //       if s.process_in_.hdr_status != PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID:
  //         s.dispatched_.exception_info.v = s.process_in_.exception_info
  //         # Copy exception info
  //         s.dispatched_.exception_info.v = s.process_in_.exception_info
  //       else:
  //         s.dispatched_.rs1.v = s.read_value[0]
  //         s.dispatched_.rs1_val.v = s.process_in_.rs1_val
  //         s.dispatched_.rs2.v = s.read_value[1]
  //         s.dispatched_.rs2_val.v = s.process_in_.rs2_val
  //         s.dispatched_.rd.v = s.process_in_.rd
  //         s.dispatched_.rd_val.v = s.process_in_.rd_val
  //         s.dispatched_.execution_data.v = s.process_in_.execution_data

  // logic for set_output()
  always @ (*) begin
    dispatched_ = 0;
    dispatched_[(74)-1:0] = process_in_[(74)-1:0];
    if ((process_in_[(2)-1:0] != PIPELINE_MSG_STATUS_VALID)) begin
      dispatched_[(142)-1:74] = process_in_[(142)-1:74];
      dispatched_[(142)-1:74] = process_in_[(142)-1:74];
    end
    else begin
      dispatched_[(139)-1:75] = read_value[0];
      dispatched_[(75)-1:74] = process_in_[(75)-1:74];
      dispatched_[(204)-1:140] = read_value[1];
      dispatched_[(140)-1:139] = process_in_[(82)-1:81];
      dispatched_[(211)-1:205] = process_in_[(95)-1:89];
      dispatched_[(205)-1:204] = process_in_[(89)-1:88];
      dispatched_[(251)-1:211] = process_in_[(135)-1:95];
    end
  end


endmodule // DispatchStage_0x3d3671bf74513fd9

//-----------------------------------------------------------------------------
// GS8LALUStage17LALUDropController_0xc628584b4321be9
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"args": ["process <C> (in_: Bits(251)) -> (accepted: Bits(1), out: Bits(146))"], "kwargs": {}}
// PyMTL: verilator_xinit = zeros
module GS8LALUStage17LALUDropController_0xc628584b4321be9
(
  input  logic [   0:0] clk,
  input  logic [ 250:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 145:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // pipeline_stage temporaries
  logic   [   0:0] pipeline_stage$check_keep;
  logic   [ 250:0] pipeline_stage$in_peek_msg;
  logic   [   0:0] pipeline_stage$clk;
  logic   [   4:0] pipeline_stage$kill_notify_msg;
  logic   [   0:0] pipeline_stage$in_peek_rdy;
  logic   [   0:0] pipeline_stage$process_accepted;
  logic   [ 145:0] pipeline_stage$check_out;
  logic   [   0:0] pipeline_stage$reset;
  logic   [ 145:0] pipeline_stage$process_out;
  logic   [   0:0] pipeline_stage$take_call;
  logic   [   0:0] pipeline_stage$process_call;
  logic   [ 145:0] pipeline_stage$check_in_;
  logic   [ 145:0] pipeline_stage$peek_msg;
  logic   [   4:0] pipeline_stage$check_msg;
  logic   [   0:0] pipeline_stage$in_take_call;
  logic   [   0:0] pipeline_stage$peek_rdy;
  logic   [ 250:0] pipeline_stage$process_in_;

  PipelineStage_0x3bdbe2fe9599a701 pipeline_stage
  (
    .check_keep       ( pipeline_stage$check_keep ),
    .in_peek_msg      ( pipeline_stage$in_peek_msg ),
    .clk              ( pipeline_stage$clk ),
    .kill_notify_msg  ( pipeline_stage$kill_notify_msg ),
    .in_peek_rdy      ( pipeline_stage$in_peek_rdy ),
    .process_accepted ( pipeline_stage$process_accepted ),
    .check_out        ( pipeline_stage$check_out ),
    .reset            ( pipeline_stage$reset ),
    .process_out      ( pipeline_stage$process_out ),
    .take_call        ( pipeline_stage$take_call ),
    .process_call     ( pipeline_stage$process_call ),
    .check_in_        ( pipeline_stage$check_in_ ),
    .peek_msg         ( pipeline_stage$peek_msg ),
    .check_msg        ( pipeline_stage$check_msg ),
    .in_take_call     ( pipeline_stage$in_take_call ),
    .peek_rdy         ( pipeline_stage$peek_rdy ),
    .process_in_      ( pipeline_stage$process_in_ )
  );

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [ 145:0] drop_controller$check_in_;
  logic   [   4:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [ 145:0] drop_controller$check_out;

  PipelineKillDropController_0x52612c5d4a64ec3 drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // stage temporaries
  logic   [   0:0] stage$process_call;
  logic   [   0:0] stage$clk;
  logic   [   0:0] stage$reset;
  logic   [ 250:0] stage$process_in_;
  logic   [   0:0] stage$process_accepted;
  logic   [ 145:0] stage$process_out;

  ALUStage_0x769b55a82b6fa607 stage
  (
    .process_call     ( stage$process_call ),
    .clk              ( stage$clk ),
    .reset            ( stage$reset ),
    .process_in_      ( stage$process_in_ ),
    .process_accepted ( stage$process_accepted ),
    .process_out      ( stage$process_out )
  );

  // signal connections
  assign drop_controller$check_in_       = pipeline_stage$check_in_;
  assign drop_controller$check_msg       = pipeline_stage$check_msg;
  assign drop_controller$clk             = clk;
  assign drop_controller$reset           = reset;
  assign in_take_call                    = pipeline_stage$in_take_call;
  assign peek_msg                        = pipeline_stage$peek_msg;
  assign peek_rdy                        = pipeline_stage$peek_rdy;
  assign pipeline_stage$check_keep       = drop_controller$check_keep;
  assign pipeline_stage$check_out        = drop_controller$check_out;
  assign pipeline_stage$clk              = clk;
  assign pipeline_stage$in_peek_msg      = in_peek_msg;
  assign pipeline_stage$in_peek_rdy      = in_peek_rdy;
  assign pipeline_stage$kill_notify_msg  = kill_notify_msg;
  assign pipeline_stage$process_accepted = stage$process_accepted;
  assign pipeline_stage$process_out      = stage$process_out;
  assign pipeline_stage$reset            = reset;
  assign pipeline_stage$take_call        = take_call;
  assign stage$clk                       = clk;
  assign stage$process_call              = pipeline_stage$process_call;
  assign stage$process_in_               = pipeline_stage$process_in_;
  assign stage$reset                     = reset;



endmodule // GS8LALUStage17LALUDropController_0xc628584b4321be9

//-----------------------------------------------------------------------------
// PipelineStage_0x3bdbe2fe9599a701
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"In": 251, "Intermediate": null, "interface": "kill_notify (msg: Bits(5)) -> (); peek <R> () -> (msg: Bits(146)); take <C> () -> ()"}
// PyMTL: verilator_xinit = zeros
module PipelineStage_0x3bdbe2fe9599a701
(
  output logic [ 145:0] check_in_,
  input  logic [   0:0] check_keep,
  output logic [   4:0] check_msg,
  input  logic [ 145:0] check_out,
  input  logic [   0:0] clk,
  input  logic [ 250:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 145:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] process_accepted,
  output logic [   0:0] process_call,
  output logic [ 250:0] process_in_,
  input  logic [ 145:0] process_out,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // logic declarations
  logic   [   0:0] output_clear;
  logic   [   0:0] input_available;


  // register declarations
  logic    [   0:0] advance;
  logic    [   0:0] taking;

  // vvm temporaries
  logic   [   0:0] vvm$check_keep;
  logic   [   0:0] vvm$clk;
  logic   [   4:0] vvm$kill_notify_msg;
  logic   [ 145:0] vvm$add_msg;
  logic   [ 145:0] vvm$check_out;
  logic   [   0:0] vvm$reset;
  logic   [   0:0] vvm$add_call;
  logic   [   0:0] vvm$take_call;
  logic   [ 145:0] vvm$check_in_;
  logic   [ 145:0] vvm$peek_msg;
  logic   [   0:0] vvm$add_rdy;
  logic   [   4:0] vvm$check_msg;
  logic   [   0:0] vvm$peek_rdy;

  ValidValueManager_0x5de589db04975131 vvm
  (
    .check_keep      ( vvm$check_keep ),
    .clk             ( vvm$clk ),
    .kill_notify_msg ( vvm$kill_notify_msg ),
    .add_msg         ( vvm$add_msg ),
    .check_out       ( vvm$check_out ),
    .reset           ( vvm$reset ),
    .add_call        ( vvm$add_call ),
    .take_call       ( vvm$take_call ),
    .check_in_       ( vvm$check_in_ ),
    .peek_msg        ( vvm$peek_msg ),
    .add_rdy         ( vvm$add_rdy ),
    .check_msg       ( vvm$check_msg ),
    .peek_rdy        ( vvm$peek_rdy )
  );

  // signal connections
  assign check_in_           = vvm$check_in_;
  assign check_msg           = vvm$check_msg;
  assign in_take_call        = taking;
  assign input_available     = in_peek_rdy;
  assign output_clear        = vvm$add_rdy;
  assign peek_msg            = vvm$peek_msg;
  assign peek_rdy            = vvm$peek_rdy;
  assign process_call        = advance;
  assign process_in_         = in_peek_msg;
  assign vvm$add_call        = taking;
  assign vvm$add_msg         = process_out;
  assign vvm$check_keep      = check_keep;
  assign vvm$check_out       = check_out;
  assign vvm$clk             = clk;
  assign vvm$kill_notify_msg = kill_notify_msg;
  assign vvm$reset           = reset;
  assign vvm$take_call       = take_call;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_taking():
  //       s.taking.v = s.advance & s.process_accepted

  // logic for handle_taking()
  always @ (*) begin
    taking = (advance&process_accepted);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_advance():
  //       s.advance.v = s.output_clear and s.input_available

  // logic for handle_advance()
  always @ (*) begin
    advance = (output_clear&&input_available);
  end


endmodule // PipelineStage_0x3bdbe2fe9599a701

//-----------------------------------------------------------------------------
// ValidValueManager_0x5de589db04975131
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"interface": "kill_notify (msg: Bits(5)) -> (); peek <R> () -> (msg: Bits(146)); take <C> () -> (); add <CR> (msg: Bits(146)) -> ()"}
// PyMTL: verilator_xinit = zeros
module ValidValueManager_0x5de589db04975131
(
  input  logic [   0:0] add_call,
  input  logic [ 145:0] add_msg,
  output logic [   0:0] add_rdy,
  output logic [ 145:0] check_in_,
  input  logic [   0:0] check_keep,
  output logic [   4:0] check_msg,
  input  logic [ 145:0] check_out,
  input  logic [   0:0] clk,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 145:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // register declarations
  logic    [   0:0] output_clear;
  logic    [   0:0] output_rdy;
  logic    [   0:0] val_reg$write_data;

  // val_reg temporaries
  logic   [   0:0] val_reg$clk;
  logic   [   0:0] val_reg$reset;
  logic   [   0:0] val_reg$read_data;

  Register_0x360ff20b8ea9d7d7 val_reg
  (
    .clk        ( val_reg$clk ),
    .write_data ( val_reg$write_data ),
    .reset      ( val_reg$reset ),
    .read_data  ( val_reg$read_data )
  );

  // out_reg temporaries
  logic   [   0:0] out_reg$clk;
  logic   [   0:0] out_reg$write_call;
  logic   [ 145:0] out_reg$write_data;
  logic   [   0:0] out_reg$reset;
  logic   [ 145:0] out_reg$read_data;

  Register_0x38751671c6f2f76 out_reg
  (
    .clk        ( out_reg$clk ),
    .write_call ( out_reg$write_call ),
    .write_data ( out_reg$write_data ),
    .reset      ( out_reg$reset ),
    .read_data  ( out_reg$read_data )
  );

  // signal connections
  assign add_rdy            = output_clear;
  assign check_in_          = out_reg$read_data;
  assign check_msg          = kill_notify_msg;
  assign out_reg$clk        = clk;
  assign out_reg$reset      = reset;
  assign out_reg$write_call = add_call;
  assign out_reg$write_data = add_msg;
  assign peek_msg           = check_out;
  assign peek_rdy           = output_rdy;
  assign val_reg$clk        = clk;
  assign val_reg$reset      = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_rdy():
  //       if s.val_reg.read_data:
  //         s.output_rdy.v = s.check_keep
  //       else:
  //         s.output_rdy.v = 0

  // logic for handle_rdy()
  always @ (*) begin
    if (val_reg$read_data) begin
      output_rdy = check_keep;
    end
    else begin
      output_rdy = 0;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_clear():
  //       s.output_clear.v = not s.output_rdy or s.take_call

  // logic for handle_clear()
  always @ (*) begin
    output_clear = (!output_rdy||take_call);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_val_reg_in():
  //       if s.add_call:
  //         s.val_reg.write_data.v = 1
  //       else:
  //         s.val_reg.write_data.v = not s.output_clear

  // logic for handle_val_reg_in()
  always @ (*) begin
    if (add_call) begin
      val_reg$write_data = 1;
    end
    else begin
      val_reg$write_data = !output_clear;
    end
  end


endmodule // ValidValueManager_0x5de589db04975131

//-----------------------------------------------------------------------------
// Register_0x38751671c6f2f76
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(146)); write <C> (data: Bits(146)) -> ()", "reset_value": null}
// PyMTL: verilator_xinit = zeros
module Register_0x38751671c6f2f76
(
  input  logic [   0:0] clk,
  output logic [ 145:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [ 145:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [ 145:0] reg_value;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (update) begin
      reg_value <= write_data;
    end
    else begin
    end
  end


endmodule // Register_0x38751671c6f2f76

//-----------------------------------------------------------------------------
// PipelineKillDropController_0x52612c5d4a64ec3
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.kill_unit {"interface": "check (msg: Bits(5), in_: Bits(146)) -> (out: Bits(146), keep: Bits(1))"}
// PyMTL: verilator_xinit = zeros
module PipelineKillDropController_0x52612c5d4a64ec3
(
  input  logic [ 145:0] check_in_,
  output logic [   0:0] check_keep,
  input  logic [   4:0] check_msg,
  output logic  [ 145:0] check_out,
  input  logic [   0:0] clk,
  input  logic [   0:0] reset
);

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [   1:0] drop_controller$check_in_;
  logic   [   4:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [   1:0] drop_controller$check_out;

  KillDropController_0xccf15b584e8c1d drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // signal connections
  assign check_keep                = drop_controller$check_keep;
  assign drop_controller$check_in_ = check_in_[73:72];
  assign drop_controller$check_msg = check_msg;
  assign drop_controller$clk       = clk;
  assign drop_controller$reset     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_out():
  //       # Set the out equal to the input and then override the branch mask
  //       s.check_out.v = s.check_in_
  //       s.check_out.hdr_branch_mask.v = s.drop_controller.check_out

  // logic for handle_out()
  always @ (*) begin
    check_out = check_in_;
    check_out[(74)-1:72] = drop_controller$check_out;
  end


endmodule // PipelineKillDropController_0x52612c5d4a64ec3

//-----------------------------------------------------------------------------
// ALUStage_0x769b55a82b6fa607
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.backend.alu {"alu_interface": "process <C> (in_: Bits(251)) -> (accepted: Bits(1), out: Bits(146))"}
// PyMTL: verilator_xinit = zeros
module ALUStage_0x769b55a82b6fa607
(
  input  logic [   0:0] clk,
  output logic [   0:0] process_accepted,
  input  logic [   0:0] process_call,
  input  logic [ 250:0] process_in_,
  output logic  [ 145:0] process_out,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [  63:0] rs1_;
  logic   [  63:0] res_;
  logic   [ 250:0] msg_;
  logic   [  63:0] rs2_;
  logic   [  63:0] imm_l20_;


  // register declarations
  logic    [  63:0] alu_$exec_src0;
  logic    [  63:0] alu_$exec_src1;
  logic    [  63:0] imm_;
  logic    [  20:0] msg_imm_;
  logic    [  31:0] res_32_;
  logic    [  63:0] res_trunc_;
  logic    [  63:0] src1_;
  logic    [  31:0] src1_32_;
  logic    [  63:0] src2_;
  logic    [  31:0] src2_32_;

  // localparam declarations
  localparam ALU_FUNC_AUIPC = 4'd10;
  localparam ALU_FUNC_LUI = 4'd9;
  localparam data_len = 64;

  // alu_ temporaries
  logic   [   0:0] alu_$exec_unsigned;
  logic   [   0:0] alu_$clk;
  logic   [   3:0] alu_$exec_func;
  logic   [   0:0] alu_$exec_call;
  logic   [   0:0] alu_$reset;
  logic   [  63:0] alu_$exec_res;
  logic   [   0:0] alu_$exec_rdy;

  ALU_0x7724efd5511f1bf4 alu_
  (
    .exec_unsigned ( alu_$exec_unsigned ),
    .clk           ( alu_$clk ),
    .exec_src1     ( alu_$exec_src1 ),
    .exec_src0     ( alu_$exec_src0 ),
    .exec_func     ( alu_$exec_func ),
    .exec_call     ( alu_$exec_call ),
    .reset         ( alu_$reset ),
    .exec_res      ( alu_$exec_res ),
    .exec_rdy      ( alu_$exec_rdy )
  );

  // op_lut_ temporaries
  logic   [   0:0] op_lut_$clk;
  logic   [   0:0] op_lut_$reset;
  logic   [   3:0] op_lut_$lookup_in_;
  logic   [   3:0] op_lut_$lookup_out;
  logic   [   0:0] op_lut_$lookup_valid;

  LookupTable_0xe1ccec17650478b op_lut_
  (
    .clk          ( op_lut_$clk ),
    .reset        ( op_lut_$reset ),
    .lookup_in_   ( op_lut_$lookup_in_ ),
    .lookup_out   ( op_lut_$lookup_out ),
    .lookup_valid ( op_lut_$lookup_valid )
  );

  // signal connections
  assign alu_$clk           = clk;
  assign alu_$exec_call     = process_call;
  assign alu_$exec_func     = op_lut_$lookup_out;
  assign alu_$exec_unsigned = msg_[241:241];
  assign alu_$reset         = reset;
  assign msg_               = process_in_;
  assign op_lut_$clk        = clk;
  assign op_lut_$lookup_in_ = msg_[239:236];
  assign op_lut_$reset      = reset;
  assign process_accepted   = 1'd1;
  assign res_               = alu_$exec_res;
  assign rs1_               = msg_[138:75];
  assign rs2_               = msg_[203:140];


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def slice32():
  //       s.src1_32_.v = s.rs1_[:32]
  //       s.src2_32_.v = s.rs2_[:32]
  //       s.res_32_.v = s.res_[:32]

  // logic for slice32()
  always @ (*) begin
    src1_32_ = rs1_[(32)-1:0];
    src2_32_ = rs2_[(32)-1:0];
    res_32_ = res_[(32)-1:0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_src_res():
  //       if s.msg_.alu_msg_op32:
  //         s.src1_.v = zext(s.src1_32_,
  //                          data_len) if s.msg_.alu_msg_unsigned else sext(
  //                              s.src1_32_, data_len)
  //         s.src2_.v = zext(s.src2_32_,
  //                          data_len) if s.msg_.alu_msg_unsigned else sext(
  //                              s.src2_32_, data_len)
  //         s.res_trunc_.v = zext(s.res_32_,
  //                               data_len) if s.msg_.alu_msg_unsigned else sext(
  //                                   s.res_32_, data_len)
  //       else:
  //         s.src1_.v = s.rs1_
  //         s.src2_.v = s.rs2_
  //         s.res_trunc_.v = s.res_
  //         if s.msg_.alu_msg_func == AluFunc.ALU_FUNC_AUIPC:
  //           s.src1_.v = s.msg_.hdr_pc
  //         elif s.msg_.alu_msg_func == AluFunc.ALU_FUNC_LUI:  # LUI is a special case
  //           s.src1_.v = 0

  // logic for set_src_res()
  always @ (*) begin
    if (msg_[(241)-1:240]) begin
      src1_ = msg_[(242)-1:241] ? { { data_len-32 { 1'b0 } }, src1_32_ } : { { data_len-32 { src1_32_[31] } }, src1_32_ };
      src2_ = msg_[(242)-1:241] ? { { data_len-32 { 1'b0 } }, src2_32_ } : { { data_len-32 { src2_32_[31] } }, src2_32_ };
      res_trunc_ = msg_[(242)-1:241] ? { { data_len-32 { 1'b0 } }, res_32_ } : { { data_len-32 { res_32_[31] } }, res_32_ };
    end
    else begin
      src1_ = rs1_;
      src2_ = rs2_;
      res_trunc_ = res_;
      if ((msg_[(240)-1:236] == ALU_FUNC_AUIPC)) begin
        src1_ = msg_[(66)-1:2];
      end
      else begin
        if ((msg_[(240)-1:236] == ALU_FUNC_LUI)) begin
          src1_ = 0;
        end
        else begin
        end
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_inputs():
  //       # PYMTL_BROKEN: sext, concat, and zext only work with wires and constants
  //       s.msg_imm_.v = s.msg_.imm
  //       s.imm_.v = sext(s.msg_imm_, data_len)
  //       if s.msg_.alu_msg_func == AluFunc.ALU_FUNC_AUIPC or s.msg_.alu_msg_func == AluFunc.ALU_FUNC_LUI:
  //         s.imm_.v = s.imm_ << 12
  //       s.alu_.exec_src0.v = s.src1_
  //       s.alu_.exec_src1.v = s.src2_ if s.msg_.rs2_val else s.imm_

  // logic for set_inputs()
  always @ (*) begin
    msg_imm_ = msg_[(233)-1:212];
    imm_ = { { data_len-21 { msg_imm_[20] } }, msg_imm_ };
    if (((msg_[(240)-1:236] == ALU_FUNC_AUIPC)||(msg_[(240)-1:236] == ALU_FUNC_LUI))) begin
      imm_ = (imm_<<12);
    end
    else begin
    end
    alu_$exec_src0 = src1_;
    alu_$exec_src1 = msg_[(140)-1:139] ? src2_ : imm_;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_process_out():
  //       s.process_out.v = 0
  //       s.process_out.hdr.v = s.msg_.hdr
  //       s.process_out.result.v = s.res_trunc_
  //       s.process_out.rd.v = s.msg_.rd
  //       s.process_out.rd_val.v = s.msg_.rd_val

  // logic for set_process_out()
  always @ (*) begin
    process_out = 0;
    process_out[(74)-1:0] = msg_[(74)-1:0];
    process_out[(146)-1:82] = res_trunc_;
    process_out[(81)-1:75] = msg_[(211)-1:205];
    process_out[(75)-1:74] = msg_[(205)-1:204];
  end


endmodule // ALUStage_0x769b55a82b6fa607

//-----------------------------------------------------------------------------
// ALU_0x7724efd5511f1bf4
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.alu {"alu_interface": "exec <CR> (src0: Bits(64), src1: Bits(64), unsigned: Bits(1), func: Bits(4)) -> (res: Bits(64))"}
// PyMTL: verilator_xinit = zeros
module ALU_0x7724efd5511f1bf4
(
  input  logic [   0:0] clk,
  input  logic [   0:0] exec_call,
  input  logic [   3:0] exec_func,
  output logic [   0:0] exec_rdy,
  output logic  [  63:0] exec_res,
  input  logic [  63:0] exec_src0,
  input  logic [  63:0] exec_src1,
  input  logic [   0:0] exec_unsigned,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   3:0] func_;
  logic   [  63:0] s1_;
  logic   [  63:0] s0_;
  logic   [   0:0] usign_;


  // register declarations
  logic    [   0:0] cmp_u_;
  logic    [  63:0] res_;
  logic    [  62:0] s0_lower_;
  logic    [   0:0] s0_up_;
  logic    [  62:0] s1_lower_;
  logic    [   0:0] s1_up_;
  logic    [   5:0] shamt_;
  logic    [ 127:0] sra_;

  // localparam declarations
  localparam ALU_ADD = 4'd0;
  localparam ALU_AND = 4'd2;
  localparam ALU_OR = 4'd3;
  localparam ALU_SLL = 4'd5;
  localparam ALU_SLT = 4'd8;
  localparam ALU_SRA = 4'd7;
  localparam ALU_SRL = 4'd6;
  localparam ALU_SUB = 4'd1;
  localparam ALU_XOR = 4'd4;
  localparam CLOG2_XLEN = 6;
  localparam TWO_XLEN = 128;
  localparam XLEN_M1 = 63;
  localparam xlen = 64;

  // signal connections
  assign exec_rdy = 1'd1;
  assign func_    = exec_func;
  assign s0_      = exec_src0;
  assign s1_      = exec_src1;
  assign usign_   = exec_unsigned;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def assign_res():
  //       s.exec_res.v = s.res_

  // logic for assign_res()
  always @ (*) begin
    exec_res = res_;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_cmp():
  //       # We flip the upper most bit if signed
  //       s.s0_up_.v = s.s0_[XLEN_M1] if s.usign_ else not s.s0_[XLEN_M1]
  //       s.s1_up_.v = s.s1_[XLEN_M1] if s.usign_ else not s.s1_[XLEN_M1]
  //       s.s0_lower_.v = s.s0_[0:XLEN_M1]
  //       s.s1_lower_.v = s.s1_[0:XLEN_M1]
  //       # Now we can concat and compare
  //       s.cmp_u_.v = concat(s.s0_up_, s.s0_lower_) < concat(s.s1_up_, s.s1_lower_)

  // logic for set_cmp()
  always @ (*) begin
    s0_up_ = usign_ ? s0_[XLEN_M1] : !s0_[XLEN_M1];
    s1_up_ = usign_ ? s1_[XLEN_M1] : !s1_[XLEN_M1];
    s0_lower_ = s0_[(XLEN_M1)-1:0];
    s1_lower_ = s1_[(XLEN_M1)-1:0];
    cmp_u_ = ({ s0_up_,s0_lower_ } < { s1_up_,s1_lower_ });
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_shamt():
  //       s.shamt_.v = s.s1_[0:CLOG2_XLEN]
  //       s.sra_.v = sext(s.s0_, TWO_XLEN) >> s.shamt_

  // logic for set_shamt()
  always @ (*) begin
    shamt_ = s1_[(CLOG2_XLEN)-1:0];
    sra_ = ({ { TWO_XLEN-64 { s0_[63] } }, s0_ }>>shamt_);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def eval_comb():
  //       s.res_.v = 0
  //       if s.exec_call:
  //         if s.func_ == ALUFunc.ALU_ADD:
  //           s.res_.v = s.s0_ + s.s1_
  //         elif s.func_ == ALUFunc.ALU_SUB:
  //           s.res_.v = s.s0_ - s.s1_
  //         elif s.func_ == ALUFunc.ALU_AND:
  //           s.res_.v = s.s0_ & s.s1_
  //         elif s.func_ == ALUFunc.ALU_OR:
  //           s.res_.v = s.s0_ | s.s1_
  //         elif s.func_ == ALUFunc.ALU_XOR:
  //           s.res_.v = s.s0_ ^ s.s1_
  //         elif s.func_ == ALUFunc.ALU_SLL:
  //           s.res_.v = s.s0_ << s.shamt_
  //         elif s.func_ == ALUFunc.ALU_SRL:
  //           s.res_.v = s.s0_ >> s.shamt_
  //         elif s.func_ == ALUFunc.ALU_SRA:
  //           s.res_.v = s.sra_[:xlen]
  //         elif s.func_ == ALUFunc.ALU_SLT:
  //           s.res_.v = zext(s.cmp_u_, xlen)

  // logic for eval_comb()
  always @ (*) begin
    res_ = 0;
    if (exec_call) begin
      if ((func_ == ALU_ADD)) begin
        res_ = (s0_+s1_);
      end
      else begin
        if ((func_ == ALU_SUB)) begin
          res_ = (s0_-s1_);
        end
        else begin
          if ((func_ == ALU_AND)) begin
            res_ = (s0_&s1_);
          end
          else begin
            if ((func_ == ALU_OR)) begin
              res_ = (s0_|s1_);
            end
            else begin
              if ((func_ == ALU_XOR)) begin
                res_ = (s0_^s1_);
              end
              else begin
                if ((func_ == ALU_SLL)) begin
                  res_ = (s0_<<shamt_);
                end
                else begin
                  if ((func_ == ALU_SRL)) begin
                    res_ = (s0_>>shamt_);
                  end
                  else begin
                    if ((func_ == ALU_SRA)) begin
                      res_ = sra_[(xlen)-1:0];
                    end
                    else begin
                      if ((func_ == ALU_SLT)) begin
                        res_ = { { xlen-1 { 1'b0 } }, cmp_u_ };
                      end
                      else begin
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    else begin
    end
  end


endmodule // ALU_0x7724efd5511f1bf4

//-----------------------------------------------------------------------------
// LookupTable_0xe1ccec17650478b
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(4)) -> (valid: Bits(1), out: Bits(4))", "mapping": {"0": "0", "1": "1", "2": "5", "3": "8", "4": "4", "5": "6", "6": "7", "7": "3", "8": "2", "9": "3", "a": "0"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0xe1ccec17650478b
(
  input  logic [   0:0] clk,
  input  logic [   3:0] lookup_in_,
  output logic [   3:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   3:0] mux$mux_default;
  logic   [   3:0] mux$mux_in_$000;
  logic   [   3:0] mux$mux_in_$001;
  logic   [   3:0] mux$mux_in_$002;
  logic   [   3:0] mux$mux_in_$003;
  logic   [   3:0] mux$mux_in_$004;
  logic   [   3:0] mux$mux_in_$005;
  logic   [   3:0] mux$mux_in_$006;
  logic   [   3:0] mux$mux_in_$007;
  logic   [   3:0] mux$mux_in_$008;
  logic   [   3:0] mux$mux_in_$009;
  logic   [   3:0] mux$mux_in_$010;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   3:0] mux$mux_select;
  logic   [   3:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x7100ff7cd1b64bc0 mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .mux_in_$003 ( mux$mux_in_$003 ),
    .mux_in_$004 ( mux$mux_in_$004 ),
    .mux_in_$005 ( mux$mux_in_$005 ),
    .mux_in_$006 ( mux$mux_in_$006 ),
    .mux_in_$007 ( mux$mux_in_$007 ),
    .mux_in_$008 ( mux$mux_in_$008 ),
    .mux_in_$009 ( mux$mux_in_$009 ),
    .mux_in_$010 ( mux$mux_in_$010 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 4'd0;
  assign mux$mux_in_$000 = 4'd0;
  assign mux$mux_in_$001 = 4'd1;
  assign mux$mux_in_$002 = 4'd5;
  assign mux$mux_in_$003 = 4'd8;
  assign mux$mux_in_$004 = 4'd4;
  assign mux$mux_in_$005 = 4'd6;
  assign mux$mux_in_$006 = 4'd7;
  assign mux$mux_in_$007 = 4'd3;
  assign mux$mux_in_$008 = 4'd2;
  assign mux$mux_in_$009 = 4'd3;
  assign mux$mux_in_$010 = 4'd0;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0xe1ccec17650478b

//-----------------------------------------------------------------------------
// CaseMux_0x7100ff7cd1b64bc0
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(4), in_: Bits(4) [11], select: Bits(4)) -> (out: Bits(4), matched: Bits(1))", "svalues": ["0", "1", "2", "3", "4", "5", "6", "7", "8", "9", "a"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x7100ff7cd1b64bc0
(
  input  logic [   0:0] clk,
  input  logic [   3:0] mux_default,
  input  logic [   3:0] mux_in_$000,
  input  logic [   3:0] mux_in_$010,
  input  logic [   3:0] mux_in_$001,
  input  logic [   3:0] mux_in_$002,
  input  logic [   3:0] mux_in_$003,
  input  logic [   3:0] mux_in_$004,
  input  logic [   3:0] mux_in_$005,
  input  logic [   3:0] mux_in_$006,
  input  logic [   3:0] mux_in_$007,
  input  logic [   3:0] mux_in_$008,
  input  logic [   3:0] mux_in_$009,
  output logic [   0:0] mux_matched,
  output logic [   3:0] mux_out,
  input  logic [   3:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   3:0] out_chain$000;
  logic   [   3:0] out_chain$001;
  logic   [   3:0] out_chain$002;
  logic   [   3:0] out_chain$003;
  logic   [   3:0] out_chain$004;
  logic   [   3:0] out_chain$005;
  logic   [   3:0] out_chain$006;
  logic   [   3:0] out_chain$007;
  logic   [   3:0] out_chain$008;
  logic   [   3:0] out_chain$009;
  logic   [   3:0] out_chain$010;
  logic   [   3:0] out_chain$011;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;
  logic   [   0:0] valid_chain$003;
  logic   [   0:0] valid_chain$004;
  logic   [   0:0] valid_chain$005;
  logic   [   0:0] valid_chain$006;
  logic   [   0:0] valid_chain$007;
  logic   [   0:0] valid_chain$008;
  logic   [   0:0] valid_chain$009;
  logic   [   0:0] valid_chain$010;
  logic   [   0:0] valid_chain$011;


  // signal connections
  assign mux_matched     = valid_chain$011;
  assign mux_out         = out_chain$011;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   3:0] mux_in_[0:10];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  assign mux_in_[  3] = mux_in_$003;
  assign mux_in_[  4] = mux_in_$004;
  assign mux_in_[  5] = mux_in_$005;
  assign mux_in_[  6] = mux_in_$006;
  assign mux_in_[  7] = mux_in_$007;
  assign mux_in_[  8] = mux_in_$008;
  assign mux_in_[  9] = mux_in_$009;
  assign mux_in_[ 10] = mux_in_$010;
  logic    [   3:0] out_chain[0:11];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  assign out_chain$003 = out_chain[  3];
  assign out_chain$004 = out_chain[  4];
  assign out_chain$005 = out_chain[  5];
  assign out_chain$006 = out_chain[  6];
  assign out_chain$007 = out_chain[  7];
  assign out_chain$008 = out_chain[  8];
  assign out_chain$009 = out_chain[  9];
  assign out_chain$010 = out_chain[ 10];
  assign out_chain$011 = out_chain[ 11];
  logic    [   0:0] valid_chain[0:11];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];
  assign valid_chain$003 = valid_chain[  3];
  assign valid_chain$004 = valid_chain[  4];
  assign valid_chain$005 = valid_chain[  5];
  assign valid_chain$006 = valid_chain[  6];
  assign valid_chain$007 = valid_chain[  7];
  assign valid_chain$008 = valid_chain[  8];
  assign valid_chain$009 = valid_chain[  9];
  assign valid_chain$010 = valid_chain[ 10];
  assign valid_chain$011 = valid_chain[ 11];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 0)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 1)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 2)) begin
      out_chain[3] = mux_in_[2];
      valid_chain[3] = 1;
    end
    else begin
      out_chain[3] = out_chain[2];
      valid_chain[3] = valid_chain[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 3)) begin
      out_chain[4] = mux_in_[3];
      valid_chain[4] = 1;
    end
    else begin
      out_chain[4] = out_chain[3];
      valid_chain[4] = valid_chain[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 4)) begin
      out_chain[5] = mux_in_[4];
      valid_chain[5] = 1;
    end
    else begin
      out_chain[5] = out_chain[4];
      valid_chain[5] = valid_chain[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 5)) begin
      out_chain[6] = mux_in_[5];
      valid_chain[6] = 1;
    end
    else begin
      out_chain[6] = out_chain[5];
      valid_chain[6] = valid_chain[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 6)) begin
      out_chain[7] = mux_in_[6];
      valid_chain[7] = 1;
    end
    else begin
      out_chain[7] = out_chain[6];
      valid_chain[7] = valid_chain[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 7)) begin
      out_chain[8] = mux_in_[7];
      valid_chain[8] = 1;
    end
    else begin
      out_chain[8] = out_chain[7];
      valid_chain[8] = valid_chain[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 8)) begin
      out_chain[9] = mux_in_[8];
      valid_chain[9] = 1;
    end
    else begin
      out_chain[9] = out_chain[8];
      valid_chain[9] = valid_chain[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 9)) begin
      out_chain[10] = mux_in_[9];
      valid_chain[10] = 1;
    end
    else begin
      out_chain[10] = out_chain[9];
      valid_chain[10] = valid_chain[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 10)) begin
      out_chain[11] = mux_in_[10];
      valid_chain[11] = 1;
    end
    else begin
      out_chain[11] = out_chain[10];
      valid_chain[11] = valid_chain[10];
    end
  end


endmodule // CaseMux_0x7100ff7cd1b64bc0

//-----------------------------------------------------------------------------
// GS11LDecodeStage28LDecodeRedirectDropController_0x15fcfedd688afdf9
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"args": ["process <C> (in_: Bits(162)) -> (accepted: Bits(1), out: Bits(190))"], "kwargs": {}}
// PyMTL: verilator_xinit = zeros
module GS11LDecodeStage28LDecodeRedirectDropController_0x15fcfedd688afdf9
(
  input  logic [   0:0] clk,
  input  logic [ 161:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   0:0] kill_notify_msg,
  output logic [ 189:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // pipeline_stage temporaries
  logic   [   0:0] pipeline_stage$check_keep;
  logic   [ 161:0] pipeline_stage$in_peek_msg;
  logic   [   0:0] pipeline_stage$clk;
  logic   [   0:0] pipeline_stage$kill_notify_msg;
  logic   [   0:0] pipeline_stage$in_peek_rdy;
  logic   [   0:0] pipeline_stage$process_accepted;
  logic   [ 189:0] pipeline_stage$check_out;
  logic   [   0:0] pipeline_stage$reset;
  logic   [ 189:0] pipeline_stage$process_out;
  logic   [   0:0] pipeline_stage$take_call;
  logic   [   0:0] pipeline_stage$process_call;
  logic   [ 189:0] pipeline_stage$check_in_;
  logic   [ 189:0] pipeline_stage$peek_msg;
  logic   [   0:0] pipeline_stage$check_msg;
  logic   [   0:0] pipeline_stage$in_take_call;
  logic   [   0:0] pipeline_stage$peek_rdy;
  logic   [ 161:0] pipeline_stage$process_in_;

  PipelineStage_0x668c1685e2c88777 pipeline_stage
  (
    .check_keep       ( pipeline_stage$check_keep ),
    .in_peek_msg      ( pipeline_stage$in_peek_msg ),
    .clk              ( pipeline_stage$clk ),
    .kill_notify_msg  ( pipeline_stage$kill_notify_msg ),
    .in_peek_rdy      ( pipeline_stage$in_peek_rdy ),
    .process_accepted ( pipeline_stage$process_accepted ),
    .check_out        ( pipeline_stage$check_out ),
    .reset            ( pipeline_stage$reset ),
    .process_out      ( pipeline_stage$process_out ),
    .take_call        ( pipeline_stage$take_call ),
    .process_call     ( pipeline_stage$process_call ),
    .check_in_        ( pipeline_stage$check_in_ ),
    .peek_msg         ( pipeline_stage$peek_msg ),
    .check_msg        ( pipeline_stage$check_msg ),
    .in_take_call     ( pipeline_stage$in_take_call ),
    .peek_rdy         ( pipeline_stage$peek_rdy ),
    .process_in_      ( pipeline_stage$process_in_ )
  );

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [ 189:0] drop_controller$check_in_;
  logic   [   0:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [ 189:0] drop_controller$check_out;

  RedirectDropController_0x530f4b732e60e820 drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // stage temporaries
  logic   [   0:0] stage$process_call;
  logic   [   0:0] stage$clk;
  logic   [   0:0] stage$reset;
  logic   [ 161:0] stage$process_in_;
  logic   [   0:0] stage$process_accepted;
  logic   [ 189:0] stage$process_out;

  DecodeStage_0x1f7a587c31394a4a stage
  (
    .process_call     ( stage$process_call ),
    .clk              ( stage$clk ),
    .reset            ( stage$reset ),
    .process_in_      ( stage$process_in_ ),
    .process_accepted ( stage$process_accepted ),
    .process_out      ( stage$process_out )
  );

  // signal connections
  assign drop_controller$check_in_       = pipeline_stage$check_in_;
  assign drop_controller$check_msg       = pipeline_stage$check_msg;
  assign drop_controller$clk             = clk;
  assign drop_controller$reset           = reset;
  assign in_take_call                    = pipeline_stage$in_take_call;
  assign peek_msg                        = pipeline_stage$peek_msg;
  assign peek_rdy                        = pipeline_stage$peek_rdy;
  assign pipeline_stage$check_keep       = drop_controller$check_keep;
  assign pipeline_stage$check_out        = drop_controller$check_out;
  assign pipeline_stage$clk              = clk;
  assign pipeline_stage$in_peek_msg      = in_peek_msg;
  assign pipeline_stage$in_peek_rdy      = in_peek_rdy;
  assign pipeline_stage$kill_notify_msg  = kill_notify_msg;
  assign pipeline_stage$process_accepted = stage$process_accepted;
  assign pipeline_stage$process_out      = stage$process_out;
  assign pipeline_stage$reset            = reset;
  assign pipeline_stage$take_call        = take_call;
  assign stage$clk                       = clk;
  assign stage$process_call              = pipeline_stage$process_call;
  assign stage$process_in_               = pipeline_stage$process_in_;
  assign stage$reset                     = reset;



endmodule // GS11LDecodeStage28LDecodeRedirectDropController_0x15fcfedd688afdf9

//-----------------------------------------------------------------------------
// PipelineStage_0x668c1685e2c88777
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"In": 162, "Intermediate": null, "interface": "kill_notify (msg: Bits(1)) -> (); peek <R> () -> (msg: Bits(190)); take <C> () -> ()"}
// PyMTL: verilator_xinit = zeros
module PipelineStage_0x668c1685e2c88777
(
  output logic [ 189:0] check_in_,
  input  logic [   0:0] check_keep,
  output logic [   0:0] check_msg,
  input  logic [ 189:0] check_out,
  input  logic [   0:0] clk,
  input  logic [ 161:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   0:0] kill_notify_msg,
  output logic [ 189:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] process_accepted,
  output logic [   0:0] process_call,
  output logic [ 161:0] process_in_,
  input  logic [ 189:0] process_out,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // logic declarations
  logic   [   0:0] output_clear;
  logic   [   0:0] input_available;


  // register declarations
  logic    [   0:0] advance;
  logic    [   0:0] taking;

  // vvm temporaries
  logic   [   0:0] vvm$check_keep;
  logic   [   0:0] vvm$clk;
  logic   [   0:0] vvm$kill_notify_msg;
  logic   [ 189:0] vvm$add_msg;
  logic   [ 189:0] vvm$check_out;
  logic   [   0:0] vvm$reset;
  logic   [   0:0] vvm$add_call;
  logic   [   0:0] vvm$take_call;
  logic   [ 189:0] vvm$check_in_;
  logic   [ 189:0] vvm$peek_msg;
  logic   [   0:0] vvm$add_rdy;
  logic   [   0:0] vvm$check_msg;
  logic   [   0:0] vvm$peek_rdy;

  ValidValueManager_0x7299a82e94b45af7 vvm
  (
    .check_keep      ( vvm$check_keep ),
    .clk             ( vvm$clk ),
    .kill_notify_msg ( vvm$kill_notify_msg ),
    .add_msg         ( vvm$add_msg ),
    .check_out       ( vvm$check_out ),
    .reset           ( vvm$reset ),
    .add_call        ( vvm$add_call ),
    .take_call       ( vvm$take_call ),
    .check_in_       ( vvm$check_in_ ),
    .peek_msg        ( vvm$peek_msg ),
    .add_rdy         ( vvm$add_rdy ),
    .check_msg       ( vvm$check_msg ),
    .peek_rdy        ( vvm$peek_rdy )
  );

  // signal connections
  assign check_in_           = vvm$check_in_;
  assign check_msg           = vvm$check_msg;
  assign in_take_call        = taking;
  assign input_available     = in_peek_rdy;
  assign output_clear        = vvm$add_rdy;
  assign peek_msg            = vvm$peek_msg;
  assign peek_rdy            = vvm$peek_rdy;
  assign process_call        = advance;
  assign process_in_         = in_peek_msg;
  assign vvm$add_call        = taking;
  assign vvm$add_msg         = process_out;
  assign vvm$check_keep      = check_keep;
  assign vvm$check_out       = check_out;
  assign vvm$clk             = clk;
  assign vvm$kill_notify_msg = kill_notify_msg;
  assign vvm$reset           = reset;
  assign vvm$take_call       = take_call;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_taking():
  //       s.taking.v = s.advance & s.process_accepted

  // logic for handle_taking()
  always @ (*) begin
    taking = (advance&process_accepted);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_advance():
  //       s.advance.v = s.output_clear and s.input_available

  // logic for handle_advance()
  always @ (*) begin
    advance = (output_clear&&input_available);
  end


endmodule // PipelineStage_0x668c1685e2c88777

//-----------------------------------------------------------------------------
// ValidValueManager_0x7299a82e94b45af7
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"interface": "kill_notify (msg: Bits(1)) -> (); peek <R> () -> (msg: Bits(190)); take <C> () -> (); add <CR> (msg: Bits(190)) -> ()"}
// PyMTL: verilator_xinit = zeros
module ValidValueManager_0x7299a82e94b45af7
(
  input  logic [   0:0] add_call,
  input  logic [ 189:0] add_msg,
  output logic [   0:0] add_rdy,
  output logic [ 189:0] check_in_,
  input  logic [   0:0] check_keep,
  output logic [   0:0] check_msg,
  input  logic [ 189:0] check_out,
  input  logic [   0:0] clk,
  input  logic [   0:0] kill_notify_msg,
  output logic [ 189:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // register declarations
  logic    [   0:0] output_clear;
  logic    [   0:0] output_rdy;
  logic    [   0:0] val_reg$write_data;

  // val_reg temporaries
  logic   [   0:0] val_reg$clk;
  logic   [   0:0] val_reg$reset;
  logic   [   0:0] val_reg$read_data;

  Register_0x360ff20b8ea9d7d7 val_reg
  (
    .clk        ( val_reg$clk ),
    .write_data ( val_reg$write_data ),
    .reset      ( val_reg$reset ),
    .read_data  ( val_reg$read_data )
  );

  // out_reg temporaries
  logic   [   0:0] out_reg$clk;
  logic   [   0:0] out_reg$write_call;
  logic   [ 189:0] out_reg$write_data;
  logic   [   0:0] out_reg$reset;
  logic   [ 189:0] out_reg$read_data;

  Register_0x14b6240d75b4640c out_reg
  (
    .clk        ( out_reg$clk ),
    .write_call ( out_reg$write_call ),
    .write_data ( out_reg$write_data ),
    .reset      ( out_reg$reset ),
    .read_data  ( out_reg$read_data )
  );

  // signal connections
  assign add_rdy            = output_clear;
  assign check_in_          = out_reg$read_data;
  assign check_msg          = kill_notify_msg;
  assign out_reg$clk        = clk;
  assign out_reg$reset      = reset;
  assign out_reg$write_call = add_call;
  assign out_reg$write_data = add_msg;
  assign peek_msg           = check_out;
  assign peek_rdy           = output_rdy;
  assign val_reg$clk        = clk;
  assign val_reg$reset      = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_rdy():
  //       if s.val_reg.read_data:
  //         s.output_rdy.v = s.check_keep
  //       else:
  //         s.output_rdy.v = 0

  // logic for handle_rdy()
  always @ (*) begin
    if (val_reg$read_data) begin
      output_rdy = check_keep;
    end
    else begin
      output_rdy = 0;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_clear():
  //       s.output_clear.v = not s.output_rdy or s.take_call

  // logic for handle_clear()
  always @ (*) begin
    output_clear = (!output_rdy||take_call);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_val_reg_in():
  //       if s.add_call:
  //         s.val_reg.write_data.v = 1
  //       else:
  //         s.val_reg.write_data.v = not s.output_clear

  // logic for handle_val_reg_in()
  always @ (*) begin
    if (add_call) begin
      val_reg$write_data = 1;
    end
    else begin
      val_reg$write_data = !output_clear;
    end
  end


endmodule // ValidValueManager_0x7299a82e94b45af7

//-----------------------------------------------------------------------------
// Register_0x14b6240d75b4640c
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(190)); write <C> (data: Bits(190)) -> ()", "reset_value": null}
// PyMTL: verilator_xinit = zeros
module Register_0x14b6240d75b4640c
(
  input  logic [   0:0] clk,
  output logic [ 189:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [ 189:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [ 189:0] reg_value;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (update) begin
      reg_value <= write_data;
    end
    else begin
    end
  end


endmodule // Register_0x14b6240d75b4640c

//-----------------------------------------------------------------------------
// RedirectDropController_0x530f4b732e60e820
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.decode {"interface": "check (msg: Bits(1), in_: Bits(190)) -> (out: Bits(190), keep: Bits(1))"}
// PyMTL: verilator_xinit = zeros
module RedirectDropController_0x530f4b732e60e820
(
  input  logic [ 189:0] check_in_,
  output logic  [   0:0] check_keep,
  input  logic [   0:0] check_msg,
  output logic [ 189:0] check_out,
  input  logic [   0:0] clk,
  input  logic [   0:0] reset
);

  // signal connections
  assign check_out = check_in_;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_check_keep():
  //       s.check_keep.v = not s.check_msg

  // logic for handle_check_keep()
  always @ (*) begin
    check_keep = !check_msg;
  end


endmodule // RedirectDropController_0x530f4b732e60e820

//-----------------------------------------------------------------------------
// DecodeStage_0x1f7a587c31394a4a
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.decode {"decode_interface": "process <C> (in_: Bits(162)) -> (accepted: Bits(1), out: Bits(190))"}
// PyMTL: verilator_xinit = zeros
module DecodeStage_0x1f7a587c31394a4a
(
  input  logic [   0:0] clk,
  output logic [   0:0] process_accepted,
  input  logic [   0:0] process_call,
  input  logic [ 161:0] process_in_,
  output logic  [ 189:0] process_out,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam ILLEGAL_INSTRUCTION = 4'd2;
  localparam PIPELINE_MSG_STATUS_EXCEPTION_RAISED = 2'd1;
  localparam PIPELINE_MSG_STATUS_VALID = 2'd0;
  localparam XLEN = 64;

  // decoder temporaries
  logic   [   0:0] decoder$clk;
  logic   [  31:0] decoder$decode_inst;
  logic   [   0:0] decoder$reset;
  logic   [   2:0] decoder$decode_imm_type;
  logic   [   0:0] decoder$decode_serialize;
  logic   [  14:0] decoder$decode_result;
  logic   [   0:0] decoder$decode_imm_val;
  logic   [   0:0] decoder$decode_rd_val;
  logic   [   0:0] decoder$decode_rs2_val;
  logic   [   2:0] decoder$decode_op_class;
  logic   [   0:0] decoder$decode_success;
  logic   [   0:0] decoder$decode_speculative;
  logic   [   0:0] decoder$decode_rs1_val;

  CD115LCD9LOpDecoder11LOp32Decoder12LOpImmDecoder14LOpImm32Decoder17LOpImmShiftDecoder19LOpImm32ShiftDecoder11LMiscDecoder10LCsrDecoder13LBranchDecoder_0x6047cbf454b06e40 decoder
  (
    .clk                ( decoder$clk ),
    .decode_inst        ( decoder$decode_inst ),
    .reset              ( decoder$reset ),
    .decode_imm_type    ( decoder$decode_imm_type ),
    .decode_serialize   ( decoder$decode_serialize ),
    .decode_result      ( decoder$decode_result ),
    .decode_imm_val     ( decoder$decode_imm_val ),
    .decode_rd_val      ( decoder$decode_rd_val ),
    .decode_rs2_val     ( decoder$decode_rs2_val ),
    .decode_op_class    ( decoder$decode_op_class ),
    .decode_success     ( decoder$decode_success ),
    .decode_speculative ( decoder$decode_speculative ),
    .decode_rs1_val     ( decoder$decode_rs1_val )
  );

  // imm_decoder temporaries
  logic   [   2:0] imm_decoder$decode_type_;
  logic   [   0:0] imm_decoder$clk;
  logic   [  31:0] imm_decoder$decode_inst;
  logic   [   0:0] imm_decoder$reset;
  logic   [  20:0] imm_decoder$decode_imm;

  ImmDecoder_0x67749655d31303e2 imm_decoder
  (
    .decode_type_ ( imm_decoder$decode_type_ ),
    .clk          ( imm_decoder$clk ),
    .decode_inst  ( imm_decoder$decode_inst ),
    .reset        ( imm_decoder$reset ),
    .decode_imm   ( imm_decoder$decode_imm )
  );

  // signal connections
  assign decoder$clk              = clk;
  assign decoder$decode_inst      = process_in_[97:66];
  assign decoder$reset            = reset;
  assign imm_decoder$clk          = clk;
  assign imm_decoder$decode_inst  = process_in_[97:66];
  assign imm_decoder$decode_type_ = decoder$decode_imm_type;
  assign imm_decoder$reset        = reset;
  assign process_accepted         = 1'd1;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode():
  //       s.process_out.v = 0
  //       s.process_out.hdr.v = s.process_in_.hdr
  //
  //       if s.process_in_.hdr_status == PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID:
  //         if s.decoder.decode_success:
  //           s.process_out.pc_succ.v = s.process_in_.pc_succ
  //
  //           s.process_out.serialize.v = s.decoder.decode_serialize
  //           s.process_out.speculative.v = s.decoder.decode_speculative
  //           s.process_out.rs1_val.v = s.decoder.decode_rs1_val
  //           s.process_out.rs1.v = s.process_in_.inst_rs1
  //           s.process_out.rs2_val.v = s.decoder.decode_rs2_val
  //           s.process_out.rs2.v = s.process_in_.inst_rs2
  //           s.process_out.rd_val.v = s.decoder.decode_rd_val
  //           s.process_out.rd.v = s.process_in_.inst_rd
  //           s.process_out.imm_val.v = s.decoder.decode_imm_val
  //           s.process_out.imm.v = s.imm_decoder.decode_imm
  //           s.process_out.op_class.v = s.decoder.decode_op_class
  //           s.process_out.pipe_msg.v = s.decoder.decode_result
  //         else:
  //           s.process_out.hdr_status.v = PipelineMsgStatus.PIPELINE_MSG_STATUS_EXCEPTION_RAISED
  //           s.process_out.exception_info_mcause.v = ExceptionCode.ILLEGAL_INSTRUCTION
  //           s.process_out.exception_info_mtval.v = zext(s.process_in_.inst, XLEN)
  //       else:
  //         s.process_out.exception_info.v = s.process_in_.exception_info

  // logic for handle_decode()
  always @ (*) begin
    process_out = 0;
    process_out[(66)-1:0] = process_in_[(66)-1:0];
    if ((process_in_[(2)-1:0] == PIPELINE_MSG_STATUS_VALID)) begin
      if (decoder$decode_success) begin
        process_out[(132)-1:68] = process_in_[(162)-1:98];
        process_out[(67)-1:66] = decoder$decode_serialize;
        process_out[(68)-1:67] = decoder$decode_speculative;
        process_out[(133)-1:132] = decoder$decode_rs1_val;
        process_out[(138)-1:133] = process_in_[(86)-1:81];
        process_out[(139)-1:138] = decoder$decode_rs2_val;
        process_out[(144)-1:139] = process_in_[(91)-1:86];
        process_out[(145)-1:144] = decoder$decode_rd_val;
        process_out[(150)-1:145] = process_in_[(78)-1:73];
        process_out[(151)-1:150] = decoder$decode_imm_val;
        process_out[(172)-1:151] = imm_decoder$decode_imm;
        process_out[(175)-1:172] = decoder$decode_op_class;
        process_out[(190)-1:175] = decoder$decode_result;
      end
      else begin
        process_out[(2)-1:0] = PIPELINE_MSG_STATUS_EXCEPTION_RAISED;
        process_out[(70)-1:66] = ILLEGAL_INSTRUCTION;
        process_out[(134)-1:70] = { { XLEN-32 { 1'b0 } }, process_in_[(98)-1:66] };
      end
    end
    else begin
      process_out[(134)-1:66] = process_in_[(134)-1:66];
    end
  end


endmodule // DecodeStage_0x1f7a587c31394a4a

//-----------------------------------------------------------------------------
// CD115LCD9LOpDecoder11LOp32Decoder12LOpImmDecoder14LOpImm32Decoder17LOpImmShiftDecoder19LOpImm32ShiftDecoder11LMiscDecoder10LCsrDecoder13LBranchDecoder_0x6047cbf454b06e40
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {}
// PyMTL: verilator_xinit = zeros
module CD115LCD9LOpDecoder11LOp32Decoder12LOpImmDecoder14LOpImm32Decoder17LOpImmShiftDecoder19LOpImm32ShiftDecoder11LMiscDecoder10LCsrDecoder13LBranchDecoder_0x6047cbf454b06e40
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // decs$000 temporaries
  logic   [   0:0] decs$000$clk;
  logic   [  31:0] decs$000$decode_inst;
  logic   [   0:0] decs$000$reset;
  logic   [   2:0] decs$000$decode_imm_type;
  logic   [   0:0] decs$000$decode_serialize;
  logic   [  14:0] decs$000$decode_result;
  logic   [   0:0] decs$000$decode_imm_val;
  logic   [   0:0] decs$000$decode_rd_val;
  logic   [   0:0] decs$000$decode_rs2_val;
  logic   [   2:0] decs$000$decode_op_class;
  logic   [   0:0] decs$000$decode_success;
  logic   [   0:0] decs$000$decode_speculative;
  logic   [   0:0] decs$000$decode_rs1_val;

  CD9LOpDecoder11LOp32Decoder12LOpImmDecoder14LOpImm32Decoder17LOpImmShiftDecoder19LOpImm32ShiftDecoder11LMiscDecoder_0x6047cbf454b06e40 decs$000
  (
    .clk                ( decs$000$clk ),
    .decode_inst        ( decs$000$decode_inst ),
    .reset              ( decs$000$reset ),
    .decode_imm_type    ( decs$000$decode_imm_type ),
    .decode_serialize   ( decs$000$decode_serialize ),
    .decode_result      ( decs$000$decode_result ),
    .decode_imm_val     ( decs$000$decode_imm_val ),
    .decode_rd_val      ( decs$000$decode_rd_val ),
    .decode_rs2_val     ( decs$000$decode_rs2_val ),
    .decode_op_class    ( decs$000$decode_op_class ),
    .decode_success     ( decs$000$decode_success ),
    .decode_speculative ( decs$000$decode_speculative ),
    .decode_rs1_val     ( decs$000$decode_rs1_val )
  );

  // decs$001 temporaries
  logic   [   0:0] decs$001$clk;
  logic   [  31:0] decs$001$decode_inst;
  logic   [   0:0] decs$001$reset;
  logic   [   2:0] decs$001$decode_imm_type;
  logic   [   0:0] decs$001$decode_serialize;
  logic   [  14:0] decs$001$decode_result;
  logic   [   0:0] decs$001$decode_imm_val;
  logic   [   0:0] decs$001$decode_rd_val;
  logic   [   0:0] decs$001$decode_rs2_val;
  logic   [   2:0] decs$001$decode_op_class;
  logic   [   0:0] decs$001$decode_success;
  logic   [   0:0] decs$001$decode_speculative;
  logic   [   0:0] decs$001$decode_rs1_val;

  CsrDecoder_0x39519b5cedf33556 decs$001
  (
    .clk                ( decs$001$clk ),
    .decode_inst        ( decs$001$decode_inst ),
    .reset              ( decs$001$reset ),
    .decode_imm_type    ( decs$001$decode_imm_type ),
    .decode_serialize   ( decs$001$decode_serialize ),
    .decode_result      ( decs$001$decode_result ),
    .decode_imm_val     ( decs$001$decode_imm_val ),
    .decode_rd_val      ( decs$001$decode_rd_val ),
    .decode_rs2_val     ( decs$001$decode_rs2_val ),
    .decode_op_class    ( decs$001$decode_op_class ),
    .decode_success     ( decs$001$decode_success ),
    .decode_speculative ( decs$001$decode_speculative ),
    .decode_rs1_val     ( decs$001$decode_rs1_val )
  );

  // decs$002 temporaries
  logic   [   0:0] decs$002$clk;
  logic   [  31:0] decs$002$decode_inst;
  logic   [   0:0] decs$002$reset;
  logic   [   2:0] decs$002$decode_imm_type;
  logic   [   0:0] decs$002$decode_serialize;
  logic   [  14:0] decs$002$decode_result;
  logic   [   0:0] decs$002$decode_imm_val;
  logic   [   0:0] decs$002$decode_rd_val;
  logic   [   0:0] decs$002$decode_rs2_val;
  logic   [   2:0] decs$002$decode_op_class;
  logic   [   0:0] decs$002$decode_success;
  logic   [   0:0] decs$002$decode_speculative;
  logic   [   0:0] decs$002$decode_rs1_val;

  GenDecoderFixed_0x30e34b165e6ab78 decs$002
  (
    .clk                ( decs$002$clk ),
    .decode_inst        ( decs$002$decode_inst ),
    .reset              ( decs$002$reset ),
    .decode_imm_type    ( decs$002$decode_imm_type ),
    .decode_serialize   ( decs$002$decode_serialize ),
    .decode_result      ( decs$002$decode_result ),
    .decode_imm_val     ( decs$002$decode_imm_val ),
    .decode_rd_val      ( decs$002$decode_rd_val ),
    .decode_rs2_val     ( decs$002$decode_rs2_val ),
    .decode_op_class    ( decs$002$decode_op_class ),
    .decode_success     ( decs$002$decode_success ),
    .decode_speculative ( decs$002$decode_speculative ),
    .decode_rs1_val     ( decs$002$decode_rs1_val )
  );

  // composite_decoder temporaries
  logic   [   0:0] composite_decoder$decode_child_serialize$000;
  logic   [   0:0] composite_decoder$decode_child_serialize$001;
  logic   [   0:0] composite_decoder$decode_child_serialize$002;
  logic   [  14:0] composite_decoder$decode_child_result$000;
  logic   [  14:0] composite_decoder$decode_child_result$001;
  logic   [  14:0] composite_decoder$decode_child_result$002;
  logic   [   0:0] composite_decoder$decode_child_imm_val$000;
  logic   [   0:0] composite_decoder$decode_child_imm_val$001;
  logic   [   0:0] composite_decoder$decode_child_imm_val$002;
  logic   [   0:0] composite_decoder$clk;
  logic   [   2:0] composite_decoder$decode_child_op_class$000;
  logic   [   2:0] composite_decoder$decode_child_op_class$001;
  logic   [   2:0] composite_decoder$decode_child_op_class$002;
  logic   [  31:0] composite_decoder$decode_inst;
  logic   [   0:0] composite_decoder$decode_child_rd_val$000;
  logic   [   0:0] composite_decoder$decode_child_rd_val$001;
  logic   [   0:0] composite_decoder$decode_child_rd_val$002;
  logic   [   0:0] composite_decoder$decode_child_speculative$000;
  logic   [   0:0] composite_decoder$decode_child_speculative$001;
  logic   [   0:0] composite_decoder$decode_child_speculative$002;
  logic   [   0:0] composite_decoder$decode_child_success$000;
  logic   [   0:0] composite_decoder$decode_child_success$001;
  logic   [   0:0] composite_decoder$decode_child_success$002;
  logic   [   0:0] composite_decoder$decode_child_rs2_val$000;
  logic   [   0:0] composite_decoder$decode_child_rs2_val$001;
  logic   [   0:0] composite_decoder$decode_child_rs2_val$002;
  logic   [   0:0] composite_decoder$reset;
  logic   [   2:0] composite_decoder$decode_child_imm_type$000;
  logic   [   2:0] composite_decoder$decode_child_imm_type$001;
  logic   [   2:0] composite_decoder$decode_child_imm_type$002;
  logic   [   0:0] composite_decoder$decode_child_rs1_val$000;
  logic   [   0:0] composite_decoder$decode_child_rs1_val$001;
  logic   [   0:0] composite_decoder$decode_child_rs1_val$002;
  logic   [   2:0] composite_decoder$decode_imm_type;
  logic   [  31:0] composite_decoder$decode_child_inst$000;
  logic   [  31:0] composite_decoder$decode_child_inst$001;
  logic   [  31:0] composite_decoder$decode_child_inst$002;
  logic   [   0:0] composite_decoder$decode_serialize;
  logic   [  14:0] composite_decoder$decode_result;
  logic   [   0:0] composite_decoder$decode_imm_val;
  logic   [   0:0] composite_decoder$decode_rd_val;
  logic   [   0:0] composite_decoder$decode_rs2_val;
  logic   [   2:0] composite_decoder$decode_op_class;
  logic   [   0:0] composite_decoder$decode_success;
  logic   [   0:0] composite_decoder$decode_speculative;
  logic   [   0:0] composite_decoder$decode_rs1_val;

  CompositeDecoder_0x2c27817f250f23b4 composite_decoder
  (
    .decode_child_serialize$000   ( composite_decoder$decode_child_serialize$000 ),
    .decode_child_serialize$001   ( composite_decoder$decode_child_serialize$001 ),
    .decode_child_serialize$002   ( composite_decoder$decode_child_serialize$002 ),
    .decode_child_result$000      ( composite_decoder$decode_child_result$000 ),
    .decode_child_result$001      ( composite_decoder$decode_child_result$001 ),
    .decode_child_result$002      ( composite_decoder$decode_child_result$002 ),
    .decode_child_imm_val$000     ( composite_decoder$decode_child_imm_val$000 ),
    .decode_child_imm_val$001     ( composite_decoder$decode_child_imm_val$001 ),
    .decode_child_imm_val$002     ( composite_decoder$decode_child_imm_val$002 ),
    .clk                          ( composite_decoder$clk ),
    .decode_child_op_class$000    ( composite_decoder$decode_child_op_class$000 ),
    .decode_child_op_class$001    ( composite_decoder$decode_child_op_class$001 ),
    .decode_child_op_class$002    ( composite_decoder$decode_child_op_class$002 ),
    .decode_inst                  ( composite_decoder$decode_inst ),
    .decode_child_rd_val$000      ( composite_decoder$decode_child_rd_val$000 ),
    .decode_child_rd_val$001      ( composite_decoder$decode_child_rd_val$001 ),
    .decode_child_rd_val$002      ( composite_decoder$decode_child_rd_val$002 ),
    .decode_child_speculative$000 ( composite_decoder$decode_child_speculative$000 ),
    .decode_child_speculative$001 ( composite_decoder$decode_child_speculative$001 ),
    .decode_child_speculative$002 ( composite_decoder$decode_child_speculative$002 ),
    .decode_child_success$000     ( composite_decoder$decode_child_success$000 ),
    .decode_child_success$001     ( composite_decoder$decode_child_success$001 ),
    .decode_child_success$002     ( composite_decoder$decode_child_success$002 ),
    .decode_child_rs2_val$000     ( composite_decoder$decode_child_rs2_val$000 ),
    .decode_child_rs2_val$001     ( composite_decoder$decode_child_rs2_val$001 ),
    .decode_child_rs2_val$002     ( composite_decoder$decode_child_rs2_val$002 ),
    .reset                        ( composite_decoder$reset ),
    .decode_child_imm_type$000    ( composite_decoder$decode_child_imm_type$000 ),
    .decode_child_imm_type$001    ( composite_decoder$decode_child_imm_type$001 ),
    .decode_child_imm_type$002    ( composite_decoder$decode_child_imm_type$002 ),
    .decode_child_rs1_val$000     ( composite_decoder$decode_child_rs1_val$000 ),
    .decode_child_rs1_val$001     ( composite_decoder$decode_child_rs1_val$001 ),
    .decode_child_rs1_val$002     ( composite_decoder$decode_child_rs1_val$002 ),
    .decode_imm_type              ( composite_decoder$decode_imm_type ),
    .decode_child_inst$000        ( composite_decoder$decode_child_inst$000 ),
    .decode_child_inst$001        ( composite_decoder$decode_child_inst$001 ),
    .decode_child_inst$002        ( composite_decoder$decode_child_inst$002 ),
    .decode_serialize             ( composite_decoder$decode_serialize ),
    .decode_result                ( composite_decoder$decode_result ),
    .decode_imm_val               ( composite_decoder$decode_imm_val ),
    .decode_rd_val                ( composite_decoder$decode_rd_val ),
    .decode_rs2_val               ( composite_decoder$decode_rs2_val ),
    .decode_op_class              ( composite_decoder$decode_op_class ),
    .decode_success               ( composite_decoder$decode_success ),
    .decode_speculative           ( composite_decoder$decode_speculative ),
    .decode_rs1_val               ( composite_decoder$decode_rs1_val )
  );

  // signal connections
  assign composite_decoder$clk                          = clk;
  assign composite_decoder$decode_child_imm_type$000    = decs$000$decode_imm_type;
  assign composite_decoder$decode_child_imm_type$001    = decs$001$decode_imm_type;
  assign composite_decoder$decode_child_imm_type$002    = decs$002$decode_imm_type;
  assign composite_decoder$decode_child_imm_val$000     = decs$000$decode_imm_val;
  assign composite_decoder$decode_child_imm_val$001     = decs$001$decode_imm_val;
  assign composite_decoder$decode_child_imm_val$002     = decs$002$decode_imm_val;
  assign composite_decoder$decode_child_op_class$000    = decs$000$decode_op_class;
  assign composite_decoder$decode_child_op_class$001    = decs$001$decode_op_class;
  assign composite_decoder$decode_child_op_class$002    = decs$002$decode_op_class;
  assign composite_decoder$decode_child_rd_val$000      = decs$000$decode_rd_val;
  assign composite_decoder$decode_child_rd_val$001      = decs$001$decode_rd_val;
  assign composite_decoder$decode_child_rd_val$002      = decs$002$decode_rd_val;
  assign composite_decoder$decode_child_result$000      = decs$000$decode_result;
  assign composite_decoder$decode_child_result$001      = decs$001$decode_result;
  assign composite_decoder$decode_child_result$002      = decs$002$decode_result;
  assign composite_decoder$decode_child_rs1_val$000     = decs$000$decode_rs1_val;
  assign composite_decoder$decode_child_rs1_val$001     = decs$001$decode_rs1_val;
  assign composite_decoder$decode_child_rs1_val$002     = decs$002$decode_rs1_val;
  assign composite_decoder$decode_child_rs2_val$000     = decs$000$decode_rs2_val;
  assign composite_decoder$decode_child_rs2_val$001     = decs$001$decode_rs2_val;
  assign composite_decoder$decode_child_rs2_val$002     = decs$002$decode_rs2_val;
  assign composite_decoder$decode_child_serialize$000   = decs$000$decode_serialize;
  assign composite_decoder$decode_child_serialize$001   = decs$001$decode_serialize;
  assign composite_decoder$decode_child_serialize$002   = decs$002$decode_serialize;
  assign composite_decoder$decode_child_speculative$000 = decs$000$decode_speculative;
  assign composite_decoder$decode_child_speculative$001 = decs$001$decode_speculative;
  assign composite_decoder$decode_child_speculative$002 = decs$002$decode_speculative;
  assign composite_decoder$decode_child_success$000     = decs$000$decode_success;
  assign composite_decoder$decode_child_success$001     = decs$001$decode_success;
  assign composite_decoder$decode_child_success$002     = decs$002$decode_success;
  assign composite_decoder$decode_inst                  = decode_inst;
  assign composite_decoder$reset                        = reset;
  assign decode_imm_type                                = composite_decoder$decode_imm_type;
  assign decode_imm_val                                 = composite_decoder$decode_imm_val;
  assign decode_op_class                                = composite_decoder$decode_op_class;
  assign decode_rd_val                                  = composite_decoder$decode_rd_val;
  assign decode_result                                  = composite_decoder$decode_result;
  assign decode_rs1_val                                 = composite_decoder$decode_rs1_val;
  assign decode_rs2_val                                 = composite_decoder$decode_rs2_val;
  assign decode_serialize                               = composite_decoder$decode_serialize;
  assign decode_speculative                             = composite_decoder$decode_speculative;
  assign decode_success                                 = composite_decoder$decode_success;
  assign decs$000$clk                                   = clk;
  assign decs$000$decode_inst                           = composite_decoder$decode_child_inst$000;
  assign decs$000$reset                                 = reset;
  assign decs$001$clk                                   = clk;
  assign decs$001$decode_inst                           = composite_decoder$decode_child_inst$001;
  assign decs$001$reset                                 = reset;
  assign decs$002$clk                                   = clk;
  assign decs$002$decode_inst                           = composite_decoder$decode_child_inst$002;
  assign decs$002$reset                                 = reset;



endmodule // CD115LCD9LOpDecoder11LOp32Decoder12LOpImmDecoder14LOpImm32Decoder17LOpImmShiftDecoder19LOpImm32ShiftDecoder11LMiscDecoder10LCsrDecoder13LBranchDecoder_0x6047cbf454b06e40

//-----------------------------------------------------------------------------
// CD9LOpDecoder11LOp32Decoder12LOpImmDecoder14LOpImm32Decoder17LOpImmShiftDecoder19LOpImm32ShiftDecoder11LMiscDecoder_0x6047cbf454b06e40
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {}
// PyMTL: verilator_xinit = zeros
module CD9LOpDecoder11LOp32Decoder12LOpImmDecoder14LOpImm32Decoder17LOpImmShiftDecoder19LOpImm32ShiftDecoder11LMiscDecoder_0x6047cbf454b06e40
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // decs$000 temporaries
  logic   [   0:0] decs$000$clk;
  logic   [  31:0] decs$000$decode_inst;
  logic   [   0:0] decs$000$reset;
  logic   [   2:0] decs$000$decode_imm_type;
  logic   [   0:0] decs$000$decode_serialize;
  logic   [  14:0] decs$000$decode_result;
  logic   [   0:0] decs$000$decode_imm_val;
  logic   [   0:0] decs$000$decode_rd_val;
  logic   [   0:0] decs$000$decode_rs2_val;
  logic   [   2:0] decs$000$decode_op_class;
  logic   [   0:0] decs$000$decode_success;
  logic   [   0:0] decs$000$decode_speculative;
  logic   [   0:0] decs$000$decode_rs1_val;

  GenDecoderFixed_0x351c7b4466e4ce87 decs$000
  (
    .clk                ( decs$000$clk ),
    .decode_inst        ( decs$000$decode_inst ),
    .reset              ( decs$000$reset ),
    .decode_imm_type    ( decs$000$decode_imm_type ),
    .decode_serialize   ( decs$000$decode_serialize ),
    .decode_result      ( decs$000$decode_result ),
    .decode_imm_val     ( decs$000$decode_imm_val ),
    .decode_rd_val      ( decs$000$decode_rd_val ),
    .decode_rs2_val     ( decs$000$decode_rs2_val ),
    .decode_op_class    ( decs$000$decode_op_class ),
    .decode_success     ( decs$000$decode_success ),
    .decode_speculative ( decs$000$decode_speculative ),
    .decode_rs1_val     ( decs$000$decode_rs1_val )
  );

  // decs$001 temporaries
  logic   [   0:0] decs$001$clk;
  logic   [  31:0] decs$001$decode_inst;
  logic   [   0:0] decs$001$reset;
  logic   [   2:0] decs$001$decode_imm_type;
  logic   [   0:0] decs$001$decode_serialize;
  logic   [  14:0] decs$001$decode_result;
  logic   [   0:0] decs$001$decode_imm_val;
  logic   [   0:0] decs$001$decode_rd_val;
  logic   [   0:0] decs$001$decode_rs2_val;
  logic   [   2:0] decs$001$decode_op_class;
  logic   [   0:0] decs$001$decode_success;
  logic   [   0:0] decs$001$decode_speculative;
  logic   [   0:0] decs$001$decode_rs1_val;

  GenDecoderFixed_0x2275b27d958d3d4e decs$001
  (
    .clk                ( decs$001$clk ),
    .decode_inst        ( decs$001$decode_inst ),
    .reset              ( decs$001$reset ),
    .decode_imm_type    ( decs$001$decode_imm_type ),
    .decode_serialize   ( decs$001$decode_serialize ),
    .decode_result      ( decs$001$decode_result ),
    .decode_imm_val     ( decs$001$decode_imm_val ),
    .decode_rd_val      ( decs$001$decode_rd_val ),
    .decode_rs2_val     ( decs$001$decode_rs2_val ),
    .decode_op_class    ( decs$001$decode_op_class ),
    .decode_success     ( decs$001$decode_success ),
    .decode_speculative ( decs$001$decode_speculative ),
    .decode_rs1_val     ( decs$001$decode_rs1_val )
  );

  // decs$002 temporaries
  logic   [   0:0] decs$002$clk;
  logic   [  31:0] decs$002$decode_inst;
  logic   [   0:0] decs$002$reset;
  logic   [   2:0] decs$002$decode_imm_type;
  logic   [   0:0] decs$002$decode_serialize;
  logic   [  14:0] decs$002$decode_result;
  logic   [   0:0] decs$002$decode_imm_val;
  logic   [   0:0] decs$002$decode_rd_val;
  logic   [   0:0] decs$002$decode_rs2_val;
  logic   [   2:0] decs$002$decode_op_class;
  logic   [   0:0] decs$002$decode_success;
  logic   [   0:0] decs$002$decode_speculative;
  logic   [   0:0] decs$002$decode_rs1_val;

  GenDecoderFixed_0x53a9336ca209e43a decs$002
  (
    .clk                ( decs$002$clk ),
    .decode_inst        ( decs$002$decode_inst ),
    .reset              ( decs$002$reset ),
    .decode_imm_type    ( decs$002$decode_imm_type ),
    .decode_serialize   ( decs$002$decode_serialize ),
    .decode_result      ( decs$002$decode_result ),
    .decode_imm_val     ( decs$002$decode_imm_val ),
    .decode_rd_val      ( decs$002$decode_rd_val ),
    .decode_rs2_val     ( decs$002$decode_rs2_val ),
    .decode_op_class    ( decs$002$decode_op_class ),
    .decode_success     ( decs$002$decode_success ),
    .decode_speculative ( decs$002$decode_speculative ),
    .decode_rs1_val     ( decs$002$decode_rs1_val )
  );

  // decs$003 temporaries
  logic   [   0:0] decs$003$clk;
  logic   [  31:0] decs$003$decode_inst;
  logic   [   0:0] decs$003$reset;
  logic   [   2:0] decs$003$decode_imm_type;
  logic   [   0:0] decs$003$decode_serialize;
  logic   [  14:0] decs$003$decode_result;
  logic   [   0:0] decs$003$decode_imm_val;
  logic   [   0:0] decs$003$decode_rd_val;
  logic   [   0:0] decs$003$decode_rs2_val;
  logic   [   2:0] decs$003$decode_op_class;
  logic   [   0:0] decs$003$decode_success;
  logic   [   0:0] decs$003$decode_speculative;
  logic   [   0:0] decs$003$decode_rs1_val;

  GenDecoderFixed_0x29e217d76d82f1af decs$003
  (
    .clk                ( decs$003$clk ),
    .decode_inst        ( decs$003$decode_inst ),
    .reset              ( decs$003$reset ),
    .decode_imm_type    ( decs$003$decode_imm_type ),
    .decode_serialize   ( decs$003$decode_serialize ),
    .decode_result      ( decs$003$decode_result ),
    .decode_imm_val     ( decs$003$decode_imm_val ),
    .decode_rd_val      ( decs$003$decode_rd_val ),
    .decode_rs2_val     ( decs$003$decode_rs2_val ),
    .decode_op_class    ( decs$003$decode_op_class ),
    .decode_success     ( decs$003$decode_success ),
    .decode_speculative ( decs$003$decode_speculative ),
    .decode_rs1_val     ( decs$003$decode_rs1_val )
  );

  // decs$004 temporaries
  logic   [   0:0] decs$004$clk;
  logic   [  31:0] decs$004$decode_inst;
  logic   [   0:0] decs$004$reset;
  logic   [   2:0] decs$004$decode_imm_type;
  logic   [   0:0] decs$004$decode_serialize;
  logic   [  14:0] decs$004$decode_result;
  logic   [   0:0] decs$004$decode_imm_val;
  logic   [   0:0] decs$004$decode_rd_val;
  logic   [   0:0] decs$004$decode_rs2_val;
  logic   [   2:0] decs$004$decode_op_class;
  logic   [   0:0] decs$004$decode_success;
  logic   [   0:0] decs$004$decode_speculative;
  logic   [   0:0] decs$004$decode_rs1_val;

  GenDecoderFixed_0x2f940af682bd257 decs$004
  (
    .clk                ( decs$004$clk ),
    .decode_inst        ( decs$004$decode_inst ),
    .reset              ( decs$004$reset ),
    .decode_imm_type    ( decs$004$decode_imm_type ),
    .decode_serialize   ( decs$004$decode_serialize ),
    .decode_result      ( decs$004$decode_result ),
    .decode_imm_val     ( decs$004$decode_imm_val ),
    .decode_rd_val      ( decs$004$decode_rd_val ),
    .decode_rs2_val     ( decs$004$decode_rs2_val ),
    .decode_op_class    ( decs$004$decode_op_class ),
    .decode_success     ( decs$004$decode_success ),
    .decode_speculative ( decs$004$decode_speculative ),
    .decode_rs1_val     ( decs$004$decode_rs1_val )
  );

  // decs$005 temporaries
  logic   [   0:0] decs$005$clk;
  logic   [  31:0] decs$005$decode_inst;
  logic   [   0:0] decs$005$reset;
  logic   [   2:0] decs$005$decode_imm_type;
  logic   [   0:0] decs$005$decode_serialize;
  logic   [  14:0] decs$005$decode_result;
  logic   [   0:0] decs$005$decode_imm_val;
  logic   [   0:0] decs$005$decode_rd_val;
  logic   [   0:0] decs$005$decode_rs2_val;
  logic   [   2:0] decs$005$decode_op_class;
  logic   [   0:0] decs$005$decode_success;
  logic   [   0:0] decs$005$decode_speculative;
  logic   [   0:0] decs$005$decode_rs1_val;

  GenDecoderFixed_0x55d6eb7561f62d2e decs$005
  (
    .clk                ( decs$005$clk ),
    .decode_inst        ( decs$005$decode_inst ),
    .reset              ( decs$005$reset ),
    .decode_imm_type    ( decs$005$decode_imm_type ),
    .decode_serialize   ( decs$005$decode_serialize ),
    .decode_result      ( decs$005$decode_result ),
    .decode_imm_val     ( decs$005$decode_imm_val ),
    .decode_rd_val      ( decs$005$decode_rd_val ),
    .decode_rs2_val     ( decs$005$decode_rs2_val ),
    .decode_op_class    ( decs$005$decode_op_class ),
    .decode_success     ( decs$005$decode_success ),
    .decode_speculative ( decs$005$decode_speculative ),
    .decode_rs1_val     ( decs$005$decode_rs1_val )
  );

  // decs$006 temporaries
  logic   [   0:0] decs$006$clk;
  logic   [  31:0] decs$006$decode_inst;
  logic   [   0:0] decs$006$reset;
  logic   [   2:0] decs$006$decode_imm_type;
  logic   [   0:0] decs$006$decode_serialize;
  logic   [  14:0] decs$006$decode_result;
  logic   [   0:0] decs$006$decode_imm_val;
  logic   [   0:0] decs$006$decode_rd_val;
  logic   [   0:0] decs$006$decode_rs2_val;
  logic   [   2:0] decs$006$decode_op_class;
  logic   [   0:0] decs$006$decode_success;
  logic   [   0:0] decs$006$decode_speculative;
  logic   [   0:0] decs$006$decode_rs1_val;

  GenDecoderFixed_0x33541dea129c9660 decs$006
  (
    .clk                ( decs$006$clk ),
    .decode_inst        ( decs$006$decode_inst ),
    .reset              ( decs$006$reset ),
    .decode_imm_type    ( decs$006$decode_imm_type ),
    .decode_serialize   ( decs$006$decode_serialize ),
    .decode_result      ( decs$006$decode_result ),
    .decode_imm_val     ( decs$006$decode_imm_val ),
    .decode_rd_val      ( decs$006$decode_rd_val ),
    .decode_rs2_val     ( decs$006$decode_rs2_val ),
    .decode_op_class    ( decs$006$decode_op_class ),
    .decode_success     ( decs$006$decode_success ),
    .decode_speculative ( decs$006$decode_speculative ),
    .decode_rs1_val     ( decs$006$decode_rs1_val )
  );

  // composite_decoder temporaries
  logic   [   0:0] composite_decoder$decode_child_serialize$000;
  logic   [   0:0] composite_decoder$decode_child_serialize$001;
  logic   [   0:0] composite_decoder$decode_child_serialize$002;
  logic   [   0:0] composite_decoder$decode_child_serialize$003;
  logic   [   0:0] composite_decoder$decode_child_serialize$004;
  logic   [   0:0] composite_decoder$decode_child_serialize$005;
  logic   [   0:0] composite_decoder$decode_child_serialize$006;
  logic   [  14:0] composite_decoder$decode_child_result$000;
  logic   [  14:0] composite_decoder$decode_child_result$001;
  logic   [  14:0] composite_decoder$decode_child_result$002;
  logic   [  14:0] composite_decoder$decode_child_result$003;
  logic   [  14:0] composite_decoder$decode_child_result$004;
  logic   [  14:0] composite_decoder$decode_child_result$005;
  logic   [  14:0] composite_decoder$decode_child_result$006;
  logic   [   0:0] composite_decoder$decode_child_imm_val$000;
  logic   [   0:0] composite_decoder$decode_child_imm_val$001;
  logic   [   0:0] composite_decoder$decode_child_imm_val$002;
  logic   [   0:0] composite_decoder$decode_child_imm_val$003;
  logic   [   0:0] composite_decoder$decode_child_imm_val$004;
  logic   [   0:0] composite_decoder$decode_child_imm_val$005;
  logic   [   0:0] composite_decoder$decode_child_imm_val$006;
  logic   [   0:0] composite_decoder$clk;
  logic   [   2:0] composite_decoder$decode_child_op_class$000;
  logic   [   2:0] composite_decoder$decode_child_op_class$001;
  logic   [   2:0] composite_decoder$decode_child_op_class$002;
  logic   [   2:0] composite_decoder$decode_child_op_class$003;
  logic   [   2:0] composite_decoder$decode_child_op_class$004;
  logic   [   2:0] composite_decoder$decode_child_op_class$005;
  logic   [   2:0] composite_decoder$decode_child_op_class$006;
  logic   [  31:0] composite_decoder$decode_inst;
  logic   [   0:0] composite_decoder$decode_child_rd_val$000;
  logic   [   0:0] composite_decoder$decode_child_rd_val$001;
  logic   [   0:0] composite_decoder$decode_child_rd_val$002;
  logic   [   0:0] composite_decoder$decode_child_rd_val$003;
  logic   [   0:0] composite_decoder$decode_child_rd_val$004;
  logic   [   0:0] composite_decoder$decode_child_rd_val$005;
  logic   [   0:0] composite_decoder$decode_child_rd_val$006;
  logic   [   0:0] composite_decoder$decode_child_speculative$000;
  logic   [   0:0] composite_decoder$decode_child_speculative$001;
  logic   [   0:0] composite_decoder$decode_child_speculative$002;
  logic   [   0:0] composite_decoder$decode_child_speculative$003;
  logic   [   0:0] composite_decoder$decode_child_speculative$004;
  logic   [   0:0] composite_decoder$decode_child_speculative$005;
  logic   [   0:0] composite_decoder$decode_child_speculative$006;
  logic   [   0:0] composite_decoder$decode_child_success$000;
  logic   [   0:0] composite_decoder$decode_child_success$001;
  logic   [   0:0] composite_decoder$decode_child_success$002;
  logic   [   0:0] composite_decoder$decode_child_success$003;
  logic   [   0:0] composite_decoder$decode_child_success$004;
  logic   [   0:0] composite_decoder$decode_child_success$005;
  logic   [   0:0] composite_decoder$decode_child_success$006;
  logic   [   0:0] composite_decoder$decode_child_rs2_val$000;
  logic   [   0:0] composite_decoder$decode_child_rs2_val$001;
  logic   [   0:0] composite_decoder$decode_child_rs2_val$002;
  logic   [   0:0] composite_decoder$decode_child_rs2_val$003;
  logic   [   0:0] composite_decoder$decode_child_rs2_val$004;
  logic   [   0:0] composite_decoder$decode_child_rs2_val$005;
  logic   [   0:0] composite_decoder$decode_child_rs2_val$006;
  logic   [   0:0] composite_decoder$reset;
  logic   [   2:0] composite_decoder$decode_child_imm_type$000;
  logic   [   2:0] composite_decoder$decode_child_imm_type$001;
  logic   [   2:0] composite_decoder$decode_child_imm_type$002;
  logic   [   2:0] composite_decoder$decode_child_imm_type$003;
  logic   [   2:0] composite_decoder$decode_child_imm_type$004;
  logic   [   2:0] composite_decoder$decode_child_imm_type$005;
  logic   [   2:0] composite_decoder$decode_child_imm_type$006;
  logic   [   0:0] composite_decoder$decode_child_rs1_val$000;
  logic   [   0:0] composite_decoder$decode_child_rs1_val$001;
  logic   [   0:0] composite_decoder$decode_child_rs1_val$002;
  logic   [   0:0] composite_decoder$decode_child_rs1_val$003;
  logic   [   0:0] composite_decoder$decode_child_rs1_val$004;
  logic   [   0:0] composite_decoder$decode_child_rs1_val$005;
  logic   [   0:0] composite_decoder$decode_child_rs1_val$006;
  logic   [   2:0] composite_decoder$decode_imm_type;
  logic   [  31:0] composite_decoder$decode_child_inst$000;
  logic   [  31:0] composite_decoder$decode_child_inst$001;
  logic   [  31:0] composite_decoder$decode_child_inst$002;
  logic   [  31:0] composite_decoder$decode_child_inst$003;
  logic   [  31:0] composite_decoder$decode_child_inst$004;
  logic   [  31:0] composite_decoder$decode_child_inst$005;
  logic   [  31:0] composite_decoder$decode_child_inst$006;
  logic   [   0:0] composite_decoder$decode_serialize;
  logic   [  14:0] composite_decoder$decode_result;
  logic   [   0:0] composite_decoder$decode_imm_val;
  logic   [   0:0] composite_decoder$decode_rd_val;
  logic   [   0:0] composite_decoder$decode_rs2_val;
  logic   [   2:0] composite_decoder$decode_op_class;
  logic   [   0:0] composite_decoder$decode_success;
  logic   [   0:0] composite_decoder$decode_speculative;
  logic   [   0:0] composite_decoder$decode_rs1_val;

  CompositeDecoder_0x2c27817f254c2cc0 composite_decoder
  (
    .decode_child_serialize$000   ( composite_decoder$decode_child_serialize$000 ),
    .decode_child_serialize$001   ( composite_decoder$decode_child_serialize$001 ),
    .decode_child_serialize$002   ( composite_decoder$decode_child_serialize$002 ),
    .decode_child_serialize$003   ( composite_decoder$decode_child_serialize$003 ),
    .decode_child_serialize$004   ( composite_decoder$decode_child_serialize$004 ),
    .decode_child_serialize$005   ( composite_decoder$decode_child_serialize$005 ),
    .decode_child_serialize$006   ( composite_decoder$decode_child_serialize$006 ),
    .decode_child_result$000      ( composite_decoder$decode_child_result$000 ),
    .decode_child_result$001      ( composite_decoder$decode_child_result$001 ),
    .decode_child_result$002      ( composite_decoder$decode_child_result$002 ),
    .decode_child_result$003      ( composite_decoder$decode_child_result$003 ),
    .decode_child_result$004      ( composite_decoder$decode_child_result$004 ),
    .decode_child_result$005      ( composite_decoder$decode_child_result$005 ),
    .decode_child_result$006      ( composite_decoder$decode_child_result$006 ),
    .decode_child_imm_val$000     ( composite_decoder$decode_child_imm_val$000 ),
    .decode_child_imm_val$001     ( composite_decoder$decode_child_imm_val$001 ),
    .decode_child_imm_val$002     ( composite_decoder$decode_child_imm_val$002 ),
    .decode_child_imm_val$003     ( composite_decoder$decode_child_imm_val$003 ),
    .decode_child_imm_val$004     ( composite_decoder$decode_child_imm_val$004 ),
    .decode_child_imm_val$005     ( composite_decoder$decode_child_imm_val$005 ),
    .decode_child_imm_val$006     ( composite_decoder$decode_child_imm_val$006 ),
    .clk                          ( composite_decoder$clk ),
    .decode_child_op_class$000    ( composite_decoder$decode_child_op_class$000 ),
    .decode_child_op_class$001    ( composite_decoder$decode_child_op_class$001 ),
    .decode_child_op_class$002    ( composite_decoder$decode_child_op_class$002 ),
    .decode_child_op_class$003    ( composite_decoder$decode_child_op_class$003 ),
    .decode_child_op_class$004    ( composite_decoder$decode_child_op_class$004 ),
    .decode_child_op_class$005    ( composite_decoder$decode_child_op_class$005 ),
    .decode_child_op_class$006    ( composite_decoder$decode_child_op_class$006 ),
    .decode_inst                  ( composite_decoder$decode_inst ),
    .decode_child_rd_val$000      ( composite_decoder$decode_child_rd_val$000 ),
    .decode_child_rd_val$001      ( composite_decoder$decode_child_rd_val$001 ),
    .decode_child_rd_val$002      ( composite_decoder$decode_child_rd_val$002 ),
    .decode_child_rd_val$003      ( composite_decoder$decode_child_rd_val$003 ),
    .decode_child_rd_val$004      ( composite_decoder$decode_child_rd_val$004 ),
    .decode_child_rd_val$005      ( composite_decoder$decode_child_rd_val$005 ),
    .decode_child_rd_val$006      ( composite_decoder$decode_child_rd_val$006 ),
    .decode_child_speculative$000 ( composite_decoder$decode_child_speculative$000 ),
    .decode_child_speculative$001 ( composite_decoder$decode_child_speculative$001 ),
    .decode_child_speculative$002 ( composite_decoder$decode_child_speculative$002 ),
    .decode_child_speculative$003 ( composite_decoder$decode_child_speculative$003 ),
    .decode_child_speculative$004 ( composite_decoder$decode_child_speculative$004 ),
    .decode_child_speculative$005 ( composite_decoder$decode_child_speculative$005 ),
    .decode_child_speculative$006 ( composite_decoder$decode_child_speculative$006 ),
    .decode_child_success$000     ( composite_decoder$decode_child_success$000 ),
    .decode_child_success$001     ( composite_decoder$decode_child_success$001 ),
    .decode_child_success$002     ( composite_decoder$decode_child_success$002 ),
    .decode_child_success$003     ( composite_decoder$decode_child_success$003 ),
    .decode_child_success$004     ( composite_decoder$decode_child_success$004 ),
    .decode_child_success$005     ( composite_decoder$decode_child_success$005 ),
    .decode_child_success$006     ( composite_decoder$decode_child_success$006 ),
    .decode_child_rs2_val$000     ( composite_decoder$decode_child_rs2_val$000 ),
    .decode_child_rs2_val$001     ( composite_decoder$decode_child_rs2_val$001 ),
    .decode_child_rs2_val$002     ( composite_decoder$decode_child_rs2_val$002 ),
    .decode_child_rs2_val$003     ( composite_decoder$decode_child_rs2_val$003 ),
    .decode_child_rs2_val$004     ( composite_decoder$decode_child_rs2_val$004 ),
    .decode_child_rs2_val$005     ( composite_decoder$decode_child_rs2_val$005 ),
    .decode_child_rs2_val$006     ( composite_decoder$decode_child_rs2_val$006 ),
    .reset                        ( composite_decoder$reset ),
    .decode_child_imm_type$000    ( composite_decoder$decode_child_imm_type$000 ),
    .decode_child_imm_type$001    ( composite_decoder$decode_child_imm_type$001 ),
    .decode_child_imm_type$002    ( composite_decoder$decode_child_imm_type$002 ),
    .decode_child_imm_type$003    ( composite_decoder$decode_child_imm_type$003 ),
    .decode_child_imm_type$004    ( composite_decoder$decode_child_imm_type$004 ),
    .decode_child_imm_type$005    ( composite_decoder$decode_child_imm_type$005 ),
    .decode_child_imm_type$006    ( composite_decoder$decode_child_imm_type$006 ),
    .decode_child_rs1_val$000     ( composite_decoder$decode_child_rs1_val$000 ),
    .decode_child_rs1_val$001     ( composite_decoder$decode_child_rs1_val$001 ),
    .decode_child_rs1_val$002     ( composite_decoder$decode_child_rs1_val$002 ),
    .decode_child_rs1_val$003     ( composite_decoder$decode_child_rs1_val$003 ),
    .decode_child_rs1_val$004     ( composite_decoder$decode_child_rs1_val$004 ),
    .decode_child_rs1_val$005     ( composite_decoder$decode_child_rs1_val$005 ),
    .decode_child_rs1_val$006     ( composite_decoder$decode_child_rs1_val$006 ),
    .decode_imm_type              ( composite_decoder$decode_imm_type ),
    .decode_child_inst$000        ( composite_decoder$decode_child_inst$000 ),
    .decode_child_inst$001        ( composite_decoder$decode_child_inst$001 ),
    .decode_child_inst$002        ( composite_decoder$decode_child_inst$002 ),
    .decode_child_inst$003        ( composite_decoder$decode_child_inst$003 ),
    .decode_child_inst$004        ( composite_decoder$decode_child_inst$004 ),
    .decode_child_inst$005        ( composite_decoder$decode_child_inst$005 ),
    .decode_child_inst$006        ( composite_decoder$decode_child_inst$006 ),
    .decode_serialize             ( composite_decoder$decode_serialize ),
    .decode_result                ( composite_decoder$decode_result ),
    .decode_imm_val               ( composite_decoder$decode_imm_val ),
    .decode_rd_val                ( composite_decoder$decode_rd_val ),
    .decode_rs2_val               ( composite_decoder$decode_rs2_val ),
    .decode_op_class              ( composite_decoder$decode_op_class ),
    .decode_success               ( composite_decoder$decode_success ),
    .decode_speculative           ( composite_decoder$decode_speculative ),
    .decode_rs1_val               ( composite_decoder$decode_rs1_val )
  );

  // signal connections
  assign composite_decoder$clk                          = clk;
  assign composite_decoder$decode_child_imm_type$000    = decs$000$decode_imm_type;
  assign composite_decoder$decode_child_imm_type$001    = decs$001$decode_imm_type;
  assign composite_decoder$decode_child_imm_type$002    = decs$002$decode_imm_type;
  assign composite_decoder$decode_child_imm_type$003    = decs$003$decode_imm_type;
  assign composite_decoder$decode_child_imm_type$004    = decs$004$decode_imm_type;
  assign composite_decoder$decode_child_imm_type$005    = decs$005$decode_imm_type;
  assign composite_decoder$decode_child_imm_type$006    = decs$006$decode_imm_type;
  assign composite_decoder$decode_child_imm_val$000     = decs$000$decode_imm_val;
  assign composite_decoder$decode_child_imm_val$001     = decs$001$decode_imm_val;
  assign composite_decoder$decode_child_imm_val$002     = decs$002$decode_imm_val;
  assign composite_decoder$decode_child_imm_val$003     = decs$003$decode_imm_val;
  assign composite_decoder$decode_child_imm_val$004     = decs$004$decode_imm_val;
  assign composite_decoder$decode_child_imm_val$005     = decs$005$decode_imm_val;
  assign composite_decoder$decode_child_imm_val$006     = decs$006$decode_imm_val;
  assign composite_decoder$decode_child_op_class$000    = decs$000$decode_op_class;
  assign composite_decoder$decode_child_op_class$001    = decs$001$decode_op_class;
  assign composite_decoder$decode_child_op_class$002    = decs$002$decode_op_class;
  assign composite_decoder$decode_child_op_class$003    = decs$003$decode_op_class;
  assign composite_decoder$decode_child_op_class$004    = decs$004$decode_op_class;
  assign composite_decoder$decode_child_op_class$005    = decs$005$decode_op_class;
  assign composite_decoder$decode_child_op_class$006    = decs$006$decode_op_class;
  assign composite_decoder$decode_child_rd_val$000      = decs$000$decode_rd_val;
  assign composite_decoder$decode_child_rd_val$001      = decs$001$decode_rd_val;
  assign composite_decoder$decode_child_rd_val$002      = decs$002$decode_rd_val;
  assign composite_decoder$decode_child_rd_val$003      = decs$003$decode_rd_val;
  assign composite_decoder$decode_child_rd_val$004      = decs$004$decode_rd_val;
  assign composite_decoder$decode_child_rd_val$005      = decs$005$decode_rd_val;
  assign composite_decoder$decode_child_rd_val$006      = decs$006$decode_rd_val;
  assign composite_decoder$decode_child_result$000      = decs$000$decode_result;
  assign composite_decoder$decode_child_result$001      = decs$001$decode_result;
  assign composite_decoder$decode_child_result$002      = decs$002$decode_result;
  assign composite_decoder$decode_child_result$003      = decs$003$decode_result;
  assign composite_decoder$decode_child_result$004      = decs$004$decode_result;
  assign composite_decoder$decode_child_result$005      = decs$005$decode_result;
  assign composite_decoder$decode_child_result$006      = decs$006$decode_result;
  assign composite_decoder$decode_child_rs1_val$000     = decs$000$decode_rs1_val;
  assign composite_decoder$decode_child_rs1_val$001     = decs$001$decode_rs1_val;
  assign composite_decoder$decode_child_rs1_val$002     = decs$002$decode_rs1_val;
  assign composite_decoder$decode_child_rs1_val$003     = decs$003$decode_rs1_val;
  assign composite_decoder$decode_child_rs1_val$004     = decs$004$decode_rs1_val;
  assign composite_decoder$decode_child_rs1_val$005     = decs$005$decode_rs1_val;
  assign composite_decoder$decode_child_rs1_val$006     = decs$006$decode_rs1_val;
  assign composite_decoder$decode_child_rs2_val$000     = decs$000$decode_rs2_val;
  assign composite_decoder$decode_child_rs2_val$001     = decs$001$decode_rs2_val;
  assign composite_decoder$decode_child_rs2_val$002     = decs$002$decode_rs2_val;
  assign composite_decoder$decode_child_rs2_val$003     = decs$003$decode_rs2_val;
  assign composite_decoder$decode_child_rs2_val$004     = decs$004$decode_rs2_val;
  assign composite_decoder$decode_child_rs2_val$005     = decs$005$decode_rs2_val;
  assign composite_decoder$decode_child_rs2_val$006     = decs$006$decode_rs2_val;
  assign composite_decoder$decode_child_serialize$000   = decs$000$decode_serialize;
  assign composite_decoder$decode_child_serialize$001   = decs$001$decode_serialize;
  assign composite_decoder$decode_child_serialize$002   = decs$002$decode_serialize;
  assign composite_decoder$decode_child_serialize$003   = decs$003$decode_serialize;
  assign composite_decoder$decode_child_serialize$004   = decs$004$decode_serialize;
  assign composite_decoder$decode_child_serialize$005   = decs$005$decode_serialize;
  assign composite_decoder$decode_child_serialize$006   = decs$006$decode_serialize;
  assign composite_decoder$decode_child_speculative$000 = decs$000$decode_speculative;
  assign composite_decoder$decode_child_speculative$001 = decs$001$decode_speculative;
  assign composite_decoder$decode_child_speculative$002 = decs$002$decode_speculative;
  assign composite_decoder$decode_child_speculative$003 = decs$003$decode_speculative;
  assign composite_decoder$decode_child_speculative$004 = decs$004$decode_speculative;
  assign composite_decoder$decode_child_speculative$005 = decs$005$decode_speculative;
  assign composite_decoder$decode_child_speculative$006 = decs$006$decode_speculative;
  assign composite_decoder$decode_child_success$000     = decs$000$decode_success;
  assign composite_decoder$decode_child_success$001     = decs$001$decode_success;
  assign composite_decoder$decode_child_success$002     = decs$002$decode_success;
  assign composite_decoder$decode_child_success$003     = decs$003$decode_success;
  assign composite_decoder$decode_child_success$004     = decs$004$decode_success;
  assign composite_decoder$decode_child_success$005     = decs$005$decode_success;
  assign composite_decoder$decode_child_success$006     = decs$006$decode_success;
  assign composite_decoder$decode_inst                  = decode_inst;
  assign composite_decoder$reset                        = reset;
  assign decode_imm_type                                = composite_decoder$decode_imm_type;
  assign decode_imm_val                                 = composite_decoder$decode_imm_val;
  assign decode_op_class                                = composite_decoder$decode_op_class;
  assign decode_rd_val                                  = composite_decoder$decode_rd_val;
  assign decode_result                                  = composite_decoder$decode_result;
  assign decode_rs1_val                                 = composite_decoder$decode_rs1_val;
  assign decode_rs2_val                                 = composite_decoder$decode_rs2_val;
  assign decode_serialize                               = composite_decoder$decode_serialize;
  assign decode_speculative                             = composite_decoder$decode_speculative;
  assign decode_success                                 = composite_decoder$decode_success;
  assign decs$000$clk                                   = clk;
  assign decs$000$decode_inst                           = composite_decoder$decode_child_inst$000;
  assign decs$000$reset                                 = reset;
  assign decs$001$clk                                   = clk;
  assign decs$001$decode_inst                           = composite_decoder$decode_child_inst$001;
  assign decs$001$reset                                 = reset;
  assign decs$002$clk                                   = clk;
  assign decs$002$decode_inst                           = composite_decoder$decode_child_inst$002;
  assign decs$002$reset                                 = reset;
  assign decs$003$clk                                   = clk;
  assign decs$003$decode_inst                           = composite_decoder$decode_child_inst$003;
  assign decs$003$reset                                 = reset;
  assign decs$004$clk                                   = clk;
  assign decs$004$decode_inst                           = composite_decoder$decode_child_inst$004;
  assign decs$004$reset                                 = reset;
  assign decs$005$clk                                   = clk;
  assign decs$005$decode_inst                           = composite_decoder$decode_child_inst$005;
  assign decs$005$reset                                 = reset;
  assign decs$006$clk                                   = clk;
  assign decs$006$decode_inst                           = composite_decoder$decode_child_inst$006;
  assign decs$006$reset                                 = reset;



endmodule // CD9LOpDecoder11LOp32Decoder12LOpImmDecoder14LOpImm32Decoder17LOpImmShiftDecoder19LOpImm32ShiftDecoder11LMiscDecoder_0x6047cbf454b06e40

//-----------------------------------------------------------------------------
// GenDecoderFixed_0x351c7b4466e4ce87
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"ResultKind": 6, "field_list": ["funct7", "funct3"], "field_map": {"(0, 0)": "func=0x0:op32=0x0:unsigned=0x0", "(0, 1)": "func=0x2:op32=0x0:unsigned=0x0", "(0, 2)": "func=0x3:op32=0x0:unsigned=0x0", "(0, 3)": "func=0x3:op32=0x0:unsigned=0x1", "(0, 4)": "func=0x4:op32=0x0:unsigned=0x0", "(0, 5)": "func=0x5:op32=0x0:unsigned=0x0", "(0, 6)": "func=0x7:op32=0x0:unsigned=0x0", "(0, 7)": "func=0x8:op32=0x0:unsigned=0x0", "(32, 0)": "func=0x1:op32=0x0:unsigned=0x0", "(32, 5)": "func=0x6:op32=0x0:unsigned=0x0"}, "fixed_map": {"opcode": "33"}, "imm_type": 0, "imm_val": 0, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 1, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoderFixed_0x351c7b4466e4ce87
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // identity_generator temporaries
  logic   [  31:0] identity_generator$gen_inst;
  logic   [   5:0] identity_generator$gen_data;
  logic   [   0:0] identity_generator$clk;
  logic   [   0:0] identity_generator$reset;
  logic   [   5:0] identity_generator$gen_payload;
  logic   [   0:0] identity_generator$gen_valid;

  IdentityPayloadGenerator_0x6a756b13525a1482 identity_generator
  (
    .gen_inst    ( identity_generator$gen_inst ),
    .gen_data    ( identity_generator$gen_data ),
    .clk         ( identity_generator$clk ),
    .reset       ( identity_generator$reset ),
    .gen_payload ( identity_generator$gen_payload ),
    .gen_valid   ( identity_generator$gen_valid )
  );

  // decoder temporaries
  logic   [   0:0] decoder$clk;
  logic   [   5:0] decoder$gen_payload;
  logic   [  31:0] decoder$decode_inst;
  logic   [   0:0] decoder$gen_valid;
  logic   [   0:0] decoder$reset;
  logic   [  31:0] decoder$gen_inst;
  logic   [   2:0] decoder$decode_imm_type;
  logic   [   5:0] decoder$gen_data;
  logic   [   0:0] decoder$decode_serialize;
  logic   [  14:0] decoder$decode_result;
  logic   [   0:0] decoder$decode_imm_val;
  logic   [   0:0] decoder$decode_rd_val;
  logic   [   0:0] decoder$decode_rs2_val;
  logic   [   2:0] decoder$decode_op_class;
  logic   [   0:0] decoder$decode_success;
  logic   [   0:0] decoder$decode_speculative;
  logic   [   0:0] decoder$decode_rs1_val;

  GenDecoder_0x13b7d6217c6defb decoder
  (
    .clk                ( decoder$clk ),
    .gen_payload        ( decoder$gen_payload ),
    .decode_inst        ( decoder$decode_inst ),
    .gen_valid          ( decoder$gen_valid ),
    .reset              ( decoder$reset ),
    .gen_inst           ( decoder$gen_inst ),
    .decode_imm_type    ( decoder$decode_imm_type ),
    .gen_data           ( decoder$gen_data ),
    .decode_serialize   ( decoder$decode_serialize ),
    .decode_result      ( decoder$decode_result ),
    .decode_imm_val     ( decoder$decode_imm_val ),
    .decode_rd_val      ( decoder$decode_rd_val ),
    .decode_rs2_val     ( decoder$decode_rs2_val ),
    .decode_op_class    ( decoder$decode_op_class ),
    .decode_success     ( decoder$decode_success ),
    .decode_speculative ( decoder$decode_speculative ),
    .decode_rs1_val     ( decoder$decode_rs1_val )
  );

  // signal connections
  assign decode_imm_type             = decoder$decode_imm_type;
  assign decode_imm_val              = decoder$decode_imm_val;
  assign decode_op_class             = decoder$decode_op_class;
  assign decode_rd_val               = decoder$decode_rd_val;
  assign decode_result               = decoder$decode_result;
  assign decode_rs1_val              = decoder$decode_rs1_val;
  assign decode_rs2_val              = decoder$decode_rs2_val;
  assign decode_serialize            = decoder$decode_serialize;
  assign decode_speculative          = decoder$decode_speculative;
  assign decode_success              = decoder$decode_success;
  assign decoder$clk                 = clk;
  assign decoder$decode_inst         = decode_inst;
  assign decoder$gen_payload         = identity_generator$gen_payload;
  assign decoder$gen_valid           = identity_generator$gen_valid;
  assign decoder$reset               = reset;
  assign identity_generator$clk      = clk;
  assign identity_generator$gen_data = decoder$gen_data;
  assign identity_generator$gen_inst = decoder$gen_inst;
  assign identity_generator$reset    = reset;



endmodule // GenDecoderFixed_0x351c7b4466e4ce87

//-----------------------------------------------------------------------------
// IdentityPayloadGenerator_0x6a756b13525a1482
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"interface": "gen (inst: Bits(32), data: Bits(6)) -> (valid: Bits(1), payload: Bits(6))"}
// PyMTL: verilator_xinit = zeros
module IdentityPayloadGenerator_0x6a756b13525a1482
(
  input  logic [   0:0] clk,
  input  logic [   5:0] gen_data,
  input  logic [  31:0] gen_inst,
  output logic [   5:0] gen_payload,
  output logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // signal connections
  assign gen_payload = gen_data;
  assign gen_valid   = 1'd1;



endmodule // IdentityPayloadGenerator_0x6a756b13525a1482

//-----------------------------------------------------------------------------
// GenDecoder_0x13b7d6217c6defb
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"In": 6, "ResultKind": 6, "field_list": ["funct7", "funct3"], "field_map": {"(0, 0)": "func=0x0:op32=0x0:unsigned=0x0", "(0, 1)": "func=0x2:op32=0x0:unsigned=0x0", "(0, 2)": "func=0x3:op32=0x0:unsigned=0x0", "(0, 3)": "func=0x3:op32=0x0:unsigned=0x1", "(0, 4)": "func=0x4:op32=0x0:unsigned=0x0", "(0, 5)": "func=0x5:op32=0x0:unsigned=0x0", "(0, 6)": "func=0x7:op32=0x0:unsigned=0x0", "(0, 7)": "func=0x8:op32=0x0:unsigned=0x0", "(32, 0)": "func=0x1:op32=0x0:unsigned=0x0", "(32, 5)": "func=0x6:op32=0x0:unsigned=0x0"}, "fixed_map": {"opcode": "33"}, "imm_type": 0, "imm_val": 0, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 1, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoder_0x13b7d6217c6defb
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic  [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic  [   0:0] decode_success,
  output logic [   5:0] gen_data,
  output logic [  31:0] gen_inst,
  input  logic [   5:0] gen_payload,
  input  logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] fixed_equals$000;
  logic   [   5:0] lookup_out;


  // lut temporaries
  logic   [   0:0] lut$clk;
  logic   [   0:0] lut$reset;
  logic   [   9:0] lut$lookup_in_;
  logic   [   5:0] lut$lookup_out;
  logic   [   0:0] lut$lookup_valid;

  LookupTable_0x87cacc5ad5b49f3 lut
  (
    .clk          ( lut$clk ),
    .reset        ( lut$reset ),
    .lookup_in_   ( lut$lookup_in_ ),
    .lookup_out   ( lut$lookup_out ),
    .lookup_valid ( lut$lookup_valid )
  );

  // equals_units$000 temporaries
  logic   [   0:0] equals_units$000$clk;
  logic   [   6:0] equals_units$000$compare_in_a;
  logic   [   6:0] equals_units$000$compare_in_b;
  logic   [   0:0] equals_units$000$reset;
  logic   [   0:0] equals_units$000$compare_out;

  Equals_0x6924ce1fe1e63d28 equals_units$000
  (
    .clk          ( equals_units$000$clk ),
    .compare_in_a ( equals_units$000$compare_in_a ),
    .compare_in_b ( equals_units$000$compare_in_b ),
    .reset        ( equals_units$000$reset ),
    .compare_out  ( equals_units$000$compare_out )
  );

  // and_unit temporaries
  logic   [   0:0] and_unit$op_in_$000;
  logic   [   0:0] and_unit$op_in_$001;
  logic   [   0:0] and_unit$clk;
  logic   [   0:0] and_unit$reset;
  logic   [   0:0] and_unit$op_out;

  And_0x8e49eae68bebab2 and_unit
  (
    .op_in_$000 ( and_unit$op_in_$000 ),
    .op_in_$001 ( and_unit$op_in_$001 ),
    .clk        ( and_unit$clk ),
    .reset      ( and_unit$reset ),
    .op_out     ( and_unit$op_out )
  );

  // signal connections
  assign and_unit$clk                  = clk;
  assign and_unit$op_in_$000           = equals_units$000$compare_out;
  assign and_unit$op_in_$001           = lut$lookup_valid;
  assign and_unit$reset                = reset;
  assign decode_imm_type               = 3'd0;
  assign decode_imm_val                = 1'd0;
  assign decode_op_class               = 3'd0;
  assign decode_rd_val                 = 1'd1;
  assign decode_rs1_val                = 1'd1;
  assign decode_rs2_val                = 1'd1;
  assign decode_serialize              = 1'd0;
  assign decode_speculative            = 1'd0;
  assign equals_units$000$clk          = clk;
  assign equals_units$000$compare_in_a = decode_inst[6:0];
  assign equals_units$000$compare_in_b = 7'd51;
  assign equals_units$000$reset        = reset;
  assign gen_data                      = lookup_out;
  assign gen_inst                      = decode_inst;
  assign lookup_out                    = lut$lookup_out;
  assign lut$clk                       = clk;
  assign lut$lookup_in_[6:0]           = decode_inst[31:25];
  assign lut$lookup_in_[9:7]           = decode_inst[14:12];
  assign lut$reset                     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_result(rs=result_field_slice.start, re=result_field_slice.stop):
  //       s.decode_result.v = 0
  //       s.decode_result[rs:re].v = s.gen_payload

  // logic for connect_result()
  always @ (*) begin
    decode_result = 0;
    decode_result[(6)-1:0] = gen_payload;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_success():
  //       s.decode_success.v = s.gen_valid & s.and_unit.op_out

  // logic for compute_success()
  always @ (*) begin
    decode_success = (gen_valid&and_unit$op_out);
  end


endmodule // GenDecoder_0x13b7d6217c6defb

//-----------------------------------------------------------------------------
// LookupTable_0x87cacc5ad5b49f3
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(10)) -> (valid: Bits(1), out: Bits(6))", "mapping": {"000": "func=0x0:op32=0x0:unsigned=0x0", "020": "func=0x1:op32=0x0:unsigned=0x0", "080": "func=0x2:op32=0x0:unsigned=0x0", "100": "func=0x3:op32=0x0:unsigned=0x0", "180": "func=0x3:op32=0x0:unsigned=0x1", "200": "func=0x4:op32=0x0:unsigned=0x0", "280": "func=0x5:op32=0x0:unsigned=0x0", "2a0": "func=0x6:op32=0x0:unsigned=0x0", "300": "func=0x7:op32=0x0:unsigned=0x0", "380": "func=0x8:op32=0x0:unsigned=0x0"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0x87cacc5ad5b49f3
(
  input  logic [   0:0] clk,
  input  logic [   9:0] lookup_in_,
  output logic [   5:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   5:0] mux$mux_default;
  logic   [   5:0] mux$mux_in_$000;
  logic   [   5:0] mux$mux_in_$001;
  logic   [   5:0] mux$mux_in_$002;
  logic   [   5:0] mux$mux_in_$003;
  logic   [   5:0] mux$mux_in_$004;
  logic   [   5:0] mux$mux_in_$005;
  logic   [   5:0] mux$mux_in_$006;
  logic   [   5:0] mux$mux_in_$007;
  logic   [   5:0] mux$mux_in_$008;
  logic   [   5:0] mux$mux_in_$009;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   9:0] mux$mux_select;
  logic   [   5:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x5243dc378d44309d mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .mux_in_$003 ( mux$mux_in_$003 ),
    .mux_in_$004 ( mux$mux_in_$004 ),
    .mux_in_$005 ( mux$mux_in_$005 ),
    .mux_in_$006 ( mux$mux_in_$006 ),
    .mux_in_$007 ( mux$mux_in_$007 ),
    .mux_in_$008 ( mux$mux_in_$008 ),
    .mux_in_$009 ( mux$mux_in_$009 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 6'd0;
  assign mux$mux_in_$000 = 6'd0;
  assign mux$mux_in_$001 = 6'd1;
  assign mux$mux_in_$002 = 6'd2;
  assign mux$mux_in_$003 = 6'd3;
  assign mux$mux_in_$004 = 6'd35;
  assign mux$mux_in_$005 = 6'd4;
  assign mux$mux_in_$006 = 6'd5;
  assign mux$mux_in_$007 = 6'd6;
  assign mux$mux_in_$008 = 6'd7;
  assign mux$mux_in_$009 = 6'd8;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0x87cacc5ad5b49f3

//-----------------------------------------------------------------------------
// CaseMux_0x5243dc378d44309d
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(6), in_: Bits(6) [10], select: Bits(10)) -> (out: Bits(6), matched: Bits(1))", "svalues": ["000", "020", "080", "100", "180", "200", "280", "2a0", "300", "380"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x5243dc378d44309d
(
  input  logic [   0:0] clk,
  input  logic [   5:0] mux_default,
  input  logic [   5:0] mux_in_$000,
  input  logic [   5:0] mux_in_$001,
  input  logic [   5:0] mux_in_$002,
  input  logic [   5:0] mux_in_$003,
  input  logic [   5:0] mux_in_$004,
  input  logic [   5:0] mux_in_$005,
  input  logic [   5:0] mux_in_$006,
  input  logic [   5:0] mux_in_$007,
  input  logic [   5:0] mux_in_$008,
  input  logic [   5:0] mux_in_$009,
  output logic [   0:0] mux_matched,
  output logic [   5:0] mux_out,
  input  logic [   9:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   5:0] out_chain$000;
  logic   [   5:0] out_chain$001;
  logic   [   5:0] out_chain$002;
  logic   [   5:0] out_chain$003;
  logic   [   5:0] out_chain$004;
  logic   [   5:0] out_chain$005;
  logic   [   5:0] out_chain$006;
  logic   [   5:0] out_chain$007;
  logic   [   5:0] out_chain$008;
  logic   [   5:0] out_chain$009;
  logic   [   5:0] out_chain$010;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;
  logic   [   0:0] valid_chain$003;
  logic   [   0:0] valid_chain$004;
  logic   [   0:0] valid_chain$005;
  logic   [   0:0] valid_chain$006;
  logic   [   0:0] valid_chain$007;
  logic   [   0:0] valid_chain$008;
  logic   [   0:0] valid_chain$009;
  logic   [   0:0] valid_chain$010;


  // signal connections
  assign mux_matched     = valid_chain$010;
  assign mux_out         = out_chain$010;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   5:0] mux_in_[0:9];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  assign mux_in_[  3] = mux_in_$003;
  assign mux_in_[  4] = mux_in_$004;
  assign mux_in_[  5] = mux_in_$005;
  assign mux_in_[  6] = mux_in_$006;
  assign mux_in_[  7] = mux_in_$007;
  assign mux_in_[  8] = mux_in_$008;
  assign mux_in_[  9] = mux_in_$009;
  logic    [   5:0] out_chain[0:10];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  assign out_chain$003 = out_chain[  3];
  assign out_chain$004 = out_chain[  4];
  assign out_chain$005 = out_chain[  5];
  assign out_chain$006 = out_chain[  6];
  assign out_chain$007 = out_chain[  7];
  assign out_chain$008 = out_chain[  8];
  assign out_chain$009 = out_chain[  9];
  assign out_chain$010 = out_chain[ 10];
  logic    [   0:0] valid_chain[0:10];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];
  assign valid_chain$003 = valid_chain[  3];
  assign valid_chain$004 = valid_chain[  4];
  assign valid_chain$005 = valid_chain[  5];
  assign valid_chain$006 = valid_chain[  6];
  assign valid_chain$007 = valid_chain[  7];
  assign valid_chain$008 = valid_chain[  8];
  assign valid_chain$009 = valid_chain[  9];
  assign valid_chain$010 = valid_chain[ 10];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 0)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 32)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 128)) begin
      out_chain[3] = mux_in_[2];
      valid_chain[3] = 1;
    end
    else begin
      out_chain[3] = out_chain[2];
      valid_chain[3] = valid_chain[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 256)) begin
      out_chain[4] = mux_in_[3];
      valid_chain[4] = 1;
    end
    else begin
      out_chain[4] = out_chain[3];
      valid_chain[4] = valid_chain[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 384)) begin
      out_chain[5] = mux_in_[4];
      valid_chain[5] = 1;
    end
    else begin
      out_chain[5] = out_chain[4];
      valid_chain[5] = valid_chain[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 512)) begin
      out_chain[6] = mux_in_[5];
      valid_chain[6] = 1;
    end
    else begin
      out_chain[6] = out_chain[5];
      valid_chain[6] = valid_chain[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 640)) begin
      out_chain[7] = mux_in_[6];
      valid_chain[7] = 1;
    end
    else begin
      out_chain[7] = out_chain[6];
      valid_chain[7] = valid_chain[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 672)) begin
      out_chain[8] = mux_in_[7];
      valid_chain[8] = 1;
    end
    else begin
      out_chain[8] = out_chain[7];
      valid_chain[8] = valid_chain[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 768)) begin
      out_chain[9] = mux_in_[8];
      valid_chain[9] = 1;
    end
    else begin
      out_chain[9] = out_chain[8];
      valid_chain[9] = valid_chain[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 896)) begin
      out_chain[10] = mux_in_[9];
      valid_chain[10] = 1;
    end
    else begin
      out_chain[10] = out_chain[9];
      valid_chain[10] = valid_chain[9];
    end
  end


endmodule // CaseMux_0x5243dc378d44309d

//-----------------------------------------------------------------------------
// Equals_0x6924ce1fe1e63d28
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.logic {"interface": "compare (in_a: Bits(7), in_b: Bits(7)) -> (out: Bits(1))"}
// PyMTL: verilator_xinit = zeros
module Equals_0x6924ce1fe1e63d28
(
  input  logic [   0:0] clk,
  input  logic [   6:0] compare_in_a,
  input  logic [   6:0] compare_in_b,
  output logic  [   0:0] compare_out,
  input  logic [   0:0] reset
);



  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute():
  //       s.compare_out.v = (s.compare_in_a == s.compare_in_b)

  // logic for compute()
  always @ (*) begin
    compare_out = (compare_in_a == compare_in_b);
  end


endmodule // Equals_0x6924ce1fe1e63d28

//-----------------------------------------------------------------------------
// And_0x8e49eae68bebab2
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.logic {"interface": "op (in_: Bits(1) [2]) -> (out: Bits(1))"}
// PyMTL: verilator_xinit = zeros
module And_0x8e49eae68bebab2
(
  input  logic [   0:0] clk,
  input  logic [   0:0] op_in_$000,
  input  logic [   0:0] op_in_$001,
  output logic [   0:0] op_out,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] partials$000;
  logic   [   0:0] partials$001;


  // signal connections
  assign op_out = partials$001;

  // array declarations
  logic   [   0:0] op_in_[0:1];
  assign op_in_[  0] = op_in_$000;
  assign op_in_[  1] = op_in_$001;
  logic    [   0:0] partials[0:1];
  assign partials$000 = partials[  0];
  assign partials$001 = partials[  1];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def initial():
  //           s.partials[0].v = s.op_in_[0]

  // logic for initial()
  always @ (*) begin
    partials[0] = op_in_[0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def next(i=i, j=i - 1):
  //           s.partials[i].v = s.op_in_[i] and s.partials[j]

  // logic for next()
  always @ (*) begin
    partials[1] = (op_in_[1]&&partials[0]);
  end


endmodule // And_0x8e49eae68bebab2

//-----------------------------------------------------------------------------
// GenDecoderFixed_0x2275b27d958d3d4e
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"ResultKind": 6, "field_list": ["funct7", "funct3"], "field_map": {"(0, 0)": "func=0x0:op32=0x1:unsigned=0x0", "(0, 1)": "func=0x2:op32=0x1:unsigned=0x0", "(0, 5)": "func=0x5:op32=0x1:unsigned=0x0", "(32, 0)": "func=0x1:op32=0x1:unsigned=0x0", "(32, 5)": "func=0x6:op32=0x1:unsigned=0x0"}, "fixed_map": {"opcode": "3b"}, "imm_type": 0, "imm_val": 0, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 1, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoderFixed_0x2275b27d958d3d4e
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // identity_generator temporaries
  logic   [  31:0] identity_generator$gen_inst;
  logic   [   5:0] identity_generator$gen_data;
  logic   [   0:0] identity_generator$clk;
  logic   [   0:0] identity_generator$reset;
  logic   [   5:0] identity_generator$gen_payload;
  logic   [   0:0] identity_generator$gen_valid;

  IdentityPayloadGenerator_0x6a756b13525a1482 identity_generator
  (
    .gen_inst    ( identity_generator$gen_inst ),
    .gen_data    ( identity_generator$gen_data ),
    .clk         ( identity_generator$clk ),
    .reset       ( identity_generator$reset ),
    .gen_payload ( identity_generator$gen_payload ),
    .gen_valid   ( identity_generator$gen_valid )
  );

  // decoder temporaries
  logic   [   0:0] decoder$clk;
  logic   [   5:0] decoder$gen_payload;
  logic   [  31:0] decoder$decode_inst;
  logic   [   0:0] decoder$gen_valid;
  logic   [   0:0] decoder$reset;
  logic   [  31:0] decoder$gen_inst;
  logic   [   2:0] decoder$decode_imm_type;
  logic   [   5:0] decoder$gen_data;
  logic   [   0:0] decoder$decode_serialize;
  logic   [  14:0] decoder$decode_result;
  logic   [   0:0] decoder$decode_imm_val;
  logic   [   0:0] decoder$decode_rd_val;
  logic   [   0:0] decoder$decode_rs2_val;
  logic   [   2:0] decoder$decode_op_class;
  logic   [   0:0] decoder$decode_success;
  logic   [   0:0] decoder$decode_speculative;
  logic   [   0:0] decoder$decode_rs1_val;

  GenDecoder_0x205f8de2c87730a2 decoder
  (
    .clk                ( decoder$clk ),
    .gen_payload        ( decoder$gen_payload ),
    .decode_inst        ( decoder$decode_inst ),
    .gen_valid          ( decoder$gen_valid ),
    .reset              ( decoder$reset ),
    .gen_inst           ( decoder$gen_inst ),
    .decode_imm_type    ( decoder$decode_imm_type ),
    .gen_data           ( decoder$gen_data ),
    .decode_serialize   ( decoder$decode_serialize ),
    .decode_result      ( decoder$decode_result ),
    .decode_imm_val     ( decoder$decode_imm_val ),
    .decode_rd_val      ( decoder$decode_rd_val ),
    .decode_rs2_val     ( decoder$decode_rs2_val ),
    .decode_op_class    ( decoder$decode_op_class ),
    .decode_success     ( decoder$decode_success ),
    .decode_speculative ( decoder$decode_speculative ),
    .decode_rs1_val     ( decoder$decode_rs1_val )
  );

  // signal connections
  assign decode_imm_type             = decoder$decode_imm_type;
  assign decode_imm_val              = decoder$decode_imm_val;
  assign decode_op_class             = decoder$decode_op_class;
  assign decode_rd_val               = decoder$decode_rd_val;
  assign decode_result               = decoder$decode_result;
  assign decode_rs1_val              = decoder$decode_rs1_val;
  assign decode_rs2_val              = decoder$decode_rs2_val;
  assign decode_serialize            = decoder$decode_serialize;
  assign decode_speculative          = decoder$decode_speculative;
  assign decode_success              = decoder$decode_success;
  assign decoder$clk                 = clk;
  assign decoder$decode_inst         = decode_inst;
  assign decoder$gen_payload         = identity_generator$gen_payload;
  assign decoder$gen_valid           = identity_generator$gen_valid;
  assign decoder$reset               = reset;
  assign identity_generator$clk      = clk;
  assign identity_generator$gen_data = decoder$gen_data;
  assign identity_generator$gen_inst = decoder$gen_inst;
  assign identity_generator$reset    = reset;



endmodule // GenDecoderFixed_0x2275b27d958d3d4e

//-----------------------------------------------------------------------------
// GenDecoder_0x205f8de2c87730a2
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"In": 6, "ResultKind": 6, "field_list": ["funct7", "funct3"], "field_map": {"(0, 0)": "func=0x0:op32=0x1:unsigned=0x0", "(0, 1)": "func=0x2:op32=0x1:unsigned=0x0", "(0, 5)": "func=0x5:op32=0x1:unsigned=0x0", "(32, 0)": "func=0x1:op32=0x1:unsigned=0x0", "(32, 5)": "func=0x6:op32=0x1:unsigned=0x0"}, "fixed_map": {"opcode": "3b"}, "imm_type": 0, "imm_val": 0, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 1, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoder_0x205f8de2c87730a2
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic  [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic  [   0:0] decode_success,
  output logic [   5:0] gen_data,
  output logic [  31:0] gen_inst,
  input  logic [   5:0] gen_payload,
  input  logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] fixed_equals$000;
  logic   [   5:0] lookup_out;


  // lut temporaries
  logic   [   0:0] lut$clk;
  logic   [   0:0] lut$reset;
  logic   [   9:0] lut$lookup_in_;
  logic   [   5:0] lut$lookup_out;
  logic   [   0:0] lut$lookup_valid;

  LookupTable_0x6327758e0f8283e3 lut
  (
    .clk          ( lut$clk ),
    .reset        ( lut$reset ),
    .lookup_in_   ( lut$lookup_in_ ),
    .lookup_out   ( lut$lookup_out ),
    .lookup_valid ( lut$lookup_valid )
  );

  // equals_units$000 temporaries
  logic   [   0:0] equals_units$000$clk;
  logic   [   6:0] equals_units$000$compare_in_a;
  logic   [   6:0] equals_units$000$compare_in_b;
  logic   [   0:0] equals_units$000$reset;
  logic   [   0:0] equals_units$000$compare_out;

  Equals_0x6924ce1fe1e63d28 equals_units$000
  (
    .clk          ( equals_units$000$clk ),
    .compare_in_a ( equals_units$000$compare_in_a ),
    .compare_in_b ( equals_units$000$compare_in_b ),
    .reset        ( equals_units$000$reset ),
    .compare_out  ( equals_units$000$compare_out )
  );

  // and_unit temporaries
  logic   [   0:0] and_unit$op_in_$000;
  logic   [   0:0] and_unit$op_in_$001;
  logic   [   0:0] and_unit$clk;
  logic   [   0:0] and_unit$reset;
  logic   [   0:0] and_unit$op_out;

  And_0x8e49eae68bebab2 and_unit
  (
    .op_in_$000 ( and_unit$op_in_$000 ),
    .op_in_$001 ( and_unit$op_in_$001 ),
    .clk        ( and_unit$clk ),
    .reset      ( and_unit$reset ),
    .op_out     ( and_unit$op_out )
  );

  // signal connections
  assign and_unit$clk                  = clk;
  assign and_unit$op_in_$000           = equals_units$000$compare_out;
  assign and_unit$op_in_$001           = lut$lookup_valid;
  assign and_unit$reset                = reset;
  assign decode_imm_type               = 3'd0;
  assign decode_imm_val                = 1'd0;
  assign decode_op_class               = 3'd0;
  assign decode_rd_val                 = 1'd1;
  assign decode_rs1_val                = 1'd1;
  assign decode_rs2_val                = 1'd1;
  assign decode_serialize              = 1'd0;
  assign decode_speculative            = 1'd0;
  assign equals_units$000$clk          = clk;
  assign equals_units$000$compare_in_a = decode_inst[6:0];
  assign equals_units$000$compare_in_b = 7'd59;
  assign equals_units$000$reset        = reset;
  assign gen_data                      = lookup_out;
  assign gen_inst                      = decode_inst;
  assign lookup_out                    = lut$lookup_out;
  assign lut$clk                       = clk;
  assign lut$lookup_in_[6:0]           = decode_inst[31:25];
  assign lut$lookup_in_[9:7]           = decode_inst[14:12];
  assign lut$reset                     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_result(rs=result_field_slice.start, re=result_field_slice.stop):
  //       s.decode_result.v = 0
  //       s.decode_result[rs:re].v = s.gen_payload

  // logic for connect_result()
  always @ (*) begin
    decode_result = 0;
    decode_result[(6)-1:0] = gen_payload;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_success():
  //       s.decode_success.v = s.gen_valid & s.and_unit.op_out

  // logic for compute_success()
  always @ (*) begin
    decode_success = (gen_valid&and_unit$op_out);
  end


endmodule // GenDecoder_0x205f8de2c87730a2

//-----------------------------------------------------------------------------
// LookupTable_0x6327758e0f8283e3
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(10)) -> (valid: Bits(1), out: Bits(6))", "mapping": {"000": "func=0x0:op32=0x1:unsigned=0x0", "020": "func=0x1:op32=0x1:unsigned=0x0", "080": "func=0x2:op32=0x1:unsigned=0x0", "280": "func=0x5:op32=0x1:unsigned=0x0", "2a0": "func=0x6:op32=0x1:unsigned=0x0"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0x6327758e0f8283e3
(
  input  logic [   0:0] clk,
  input  logic [   9:0] lookup_in_,
  output logic [   5:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   5:0] mux$mux_default;
  logic   [   5:0] mux$mux_in_$000;
  logic   [   5:0] mux$mux_in_$001;
  logic   [   5:0] mux$mux_in_$002;
  logic   [   5:0] mux$mux_in_$003;
  logic   [   5:0] mux$mux_in_$004;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   9:0] mux$mux_select;
  logic   [   5:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x561022ff67649b35 mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .mux_in_$003 ( mux$mux_in_$003 ),
    .mux_in_$004 ( mux$mux_in_$004 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 6'd0;
  assign mux$mux_in_$000 = 6'd16;
  assign mux$mux_in_$001 = 6'd17;
  assign mux$mux_in_$002 = 6'd18;
  assign mux$mux_in_$003 = 6'd21;
  assign mux$mux_in_$004 = 6'd22;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0x6327758e0f8283e3

//-----------------------------------------------------------------------------
// CaseMux_0x561022ff67649b35
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(6), in_: Bits(6) [5], select: Bits(10)) -> (out: Bits(6), matched: Bits(1))", "svalues": ["000", "020", "080", "280", "2a0"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x561022ff67649b35
(
  input  logic [   0:0] clk,
  input  logic [   5:0] mux_default,
  input  logic [   5:0] mux_in_$000,
  input  logic [   5:0] mux_in_$001,
  input  logic [   5:0] mux_in_$002,
  input  logic [   5:0] mux_in_$003,
  input  logic [   5:0] mux_in_$004,
  output logic [   0:0] mux_matched,
  output logic [   5:0] mux_out,
  input  logic [   9:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   5:0] out_chain$000;
  logic   [   5:0] out_chain$001;
  logic   [   5:0] out_chain$002;
  logic   [   5:0] out_chain$003;
  logic   [   5:0] out_chain$004;
  logic   [   5:0] out_chain$005;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;
  logic   [   0:0] valid_chain$003;
  logic   [   0:0] valid_chain$004;
  logic   [   0:0] valid_chain$005;


  // signal connections
  assign mux_matched     = valid_chain$005;
  assign mux_out         = out_chain$005;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   5:0] mux_in_[0:4];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  assign mux_in_[  3] = mux_in_$003;
  assign mux_in_[  4] = mux_in_$004;
  logic    [   5:0] out_chain[0:5];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  assign out_chain$003 = out_chain[  3];
  assign out_chain$004 = out_chain[  4];
  assign out_chain$005 = out_chain[  5];
  logic    [   0:0] valid_chain[0:5];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];
  assign valid_chain$003 = valid_chain[  3];
  assign valid_chain$004 = valid_chain[  4];
  assign valid_chain$005 = valid_chain[  5];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 0)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 32)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 128)) begin
      out_chain[3] = mux_in_[2];
      valid_chain[3] = 1;
    end
    else begin
      out_chain[3] = out_chain[2];
      valid_chain[3] = valid_chain[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 640)) begin
      out_chain[4] = mux_in_[3];
      valid_chain[4] = 1;
    end
    else begin
      out_chain[4] = out_chain[3];
      valid_chain[4] = valid_chain[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 672)) begin
      out_chain[5] = mux_in_[4];
      valid_chain[5] = 1;
    end
    else begin
      out_chain[5] = out_chain[4];
      valid_chain[5] = valid_chain[4];
    end
  end


endmodule // CaseMux_0x561022ff67649b35

//-----------------------------------------------------------------------------
// GenDecoderFixed_0x53a9336ca209e43a
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"ResultKind": 6, "field_list": ["funct3"], "field_map": {"0": "func=0x0:op32=0x0:unsigned=0x0", "2": "func=0x3:op32=0x0:unsigned=0x0", "3": "func=0x3:op32=0x0:unsigned=0x1", "4": "func=0x4:op32=0x0:unsigned=0x0", "6": "func=0x7:op32=0x0:unsigned=0x0", "7": "func=0x8:op32=0x0:unsigned=0x0"}, "fixed_map": {"opcode": "13"}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 0, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoderFixed_0x53a9336ca209e43a
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // identity_generator temporaries
  logic   [  31:0] identity_generator$gen_inst;
  logic   [   5:0] identity_generator$gen_data;
  logic   [   0:0] identity_generator$clk;
  logic   [   0:0] identity_generator$reset;
  logic   [   5:0] identity_generator$gen_payload;
  logic   [   0:0] identity_generator$gen_valid;

  IdentityPayloadGenerator_0x6a756b13525a1482 identity_generator
  (
    .gen_inst    ( identity_generator$gen_inst ),
    .gen_data    ( identity_generator$gen_data ),
    .clk         ( identity_generator$clk ),
    .reset       ( identity_generator$reset ),
    .gen_payload ( identity_generator$gen_payload ),
    .gen_valid   ( identity_generator$gen_valid )
  );

  // decoder temporaries
  logic   [   0:0] decoder$clk;
  logic   [   5:0] decoder$gen_payload;
  logic   [  31:0] decoder$decode_inst;
  logic   [   0:0] decoder$gen_valid;
  logic   [   0:0] decoder$reset;
  logic   [  31:0] decoder$gen_inst;
  logic   [   2:0] decoder$decode_imm_type;
  logic   [   5:0] decoder$gen_data;
  logic   [   0:0] decoder$decode_serialize;
  logic   [  14:0] decoder$decode_result;
  logic   [   0:0] decoder$decode_imm_val;
  logic   [   0:0] decoder$decode_rd_val;
  logic   [   0:0] decoder$decode_rs2_val;
  logic   [   2:0] decoder$decode_op_class;
  logic   [   0:0] decoder$decode_success;
  logic   [   0:0] decoder$decode_speculative;
  logic   [   0:0] decoder$decode_rs1_val;

  GenDecoder_0x7d917d4fc7f6270a decoder
  (
    .clk                ( decoder$clk ),
    .gen_payload        ( decoder$gen_payload ),
    .decode_inst        ( decoder$decode_inst ),
    .gen_valid          ( decoder$gen_valid ),
    .reset              ( decoder$reset ),
    .gen_inst           ( decoder$gen_inst ),
    .decode_imm_type    ( decoder$decode_imm_type ),
    .gen_data           ( decoder$gen_data ),
    .decode_serialize   ( decoder$decode_serialize ),
    .decode_result      ( decoder$decode_result ),
    .decode_imm_val     ( decoder$decode_imm_val ),
    .decode_rd_val      ( decoder$decode_rd_val ),
    .decode_rs2_val     ( decoder$decode_rs2_val ),
    .decode_op_class    ( decoder$decode_op_class ),
    .decode_success     ( decoder$decode_success ),
    .decode_speculative ( decoder$decode_speculative ),
    .decode_rs1_val     ( decoder$decode_rs1_val )
  );

  // signal connections
  assign decode_imm_type             = decoder$decode_imm_type;
  assign decode_imm_val              = decoder$decode_imm_val;
  assign decode_op_class             = decoder$decode_op_class;
  assign decode_rd_val               = decoder$decode_rd_val;
  assign decode_result               = decoder$decode_result;
  assign decode_rs1_val              = decoder$decode_rs1_val;
  assign decode_rs2_val              = decoder$decode_rs2_val;
  assign decode_serialize            = decoder$decode_serialize;
  assign decode_speculative          = decoder$decode_speculative;
  assign decode_success              = decoder$decode_success;
  assign decoder$clk                 = clk;
  assign decoder$decode_inst         = decode_inst;
  assign decoder$gen_payload         = identity_generator$gen_payload;
  assign decoder$gen_valid           = identity_generator$gen_valid;
  assign decoder$reset               = reset;
  assign identity_generator$clk      = clk;
  assign identity_generator$gen_data = decoder$gen_data;
  assign identity_generator$gen_inst = decoder$gen_inst;
  assign identity_generator$reset    = reset;



endmodule // GenDecoderFixed_0x53a9336ca209e43a

//-----------------------------------------------------------------------------
// GenDecoder_0x7d917d4fc7f6270a
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"In": 6, "ResultKind": 6, "field_list": ["funct3"], "field_map": {"0": "func=0x0:op32=0x0:unsigned=0x0", "2": "func=0x3:op32=0x0:unsigned=0x0", "3": "func=0x3:op32=0x0:unsigned=0x1", "4": "func=0x4:op32=0x0:unsigned=0x0", "6": "func=0x7:op32=0x0:unsigned=0x0", "7": "func=0x8:op32=0x0:unsigned=0x0"}, "fixed_map": {"opcode": "13"}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 0, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoder_0x7d917d4fc7f6270a
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic  [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic  [   0:0] decode_success,
  output logic [   5:0] gen_data,
  output logic [  31:0] gen_inst,
  input  logic [   5:0] gen_payload,
  input  logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] fixed_equals$000;
  logic   [   5:0] lookup_out;


  // lut temporaries
  logic   [   0:0] lut$clk;
  logic   [   0:0] lut$reset;
  logic   [   2:0] lut$lookup_in_;
  logic   [   5:0] lut$lookup_out;
  logic   [   0:0] lut$lookup_valid;

  LookupTable_0x3f37677ed10fc59b lut
  (
    .clk          ( lut$clk ),
    .reset        ( lut$reset ),
    .lookup_in_   ( lut$lookup_in_ ),
    .lookup_out   ( lut$lookup_out ),
    .lookup_valid ( lut$lookup_valid )
  );

  // equals_units$000 temporaries
  logic   [   0:0] equals_units$000$clk;
  logic   [   6:0] equals_units$000$compare_in_a;
  logic   [   6:0] equals_units$000$compare_in_b;
  logic   [   0:0] equals_units$000$reset;
  logic   [   0:0] equals_units$000$compare_out;

  Equals_0x6924ce1fe1e63d28 equals_units$000
  (
    .clk          ( equals_units$000$clk ),
    .compare_in_a ( equals_units$000$compare_in_a ),
    .compare_in_b ( equals_units$000$compare_in_b ),
    .reset        ( equals_units$000$reset ),
    .compare_out  ( equals_units$000$compare_out )
  );

  // and_unit temporaries
  logic   [   0:0] and_unit$op_in_$000;
  logic   [   0:0] and_unit$op_in_$001;
  logic   [   0:0] and_unit$clk;
  logic   [   0:0] and_unit$reset;
  logic   [   0:0] and_unit$op_out;

  And_0x8e49eae68bebab2 and_unit
  (
    .op_in_$000 ( and_unit$op_in_$000 ),
    .op_in_$001 ( and_unit$op_in_$001 ),
    .clk        ( and_unit$clk ),
    .reset      ( and_unit$reset ),
    .op_out     ( and_unit$op_out )
  );

  // signal connections
  assign and_unit$clk                  = clk;
  assign and_unit$op_in_$000           = equals_units$000$compare_out;
  assign and_unit$op_in_$001           = lut$lookup_valid;
  assign and_unit$reset                = reset;
  assign decode_imm_type               = 3'd0;
  assign decode_imm_val                = 1'd1;
  assign decode_op_class               = 3'd0;
  assign decode_rd_val                 = 1'd1;
  assign decode_rs1_val                = 1'd1;
  assign decode_rs2_val                = 1'd0;
  assign decode_serialize              = 1'd0;
  assign decode_speculative            = 1'd0;
  assign equals_units$000$clk          = clk;
  assign equals_units$000$compare_in_a = decode_inst[6:0];
  assign equals_units$000$compare_in_b = 7'd19;
  assign equals_units$000$reset        = reset;
  assign gen_data                      = lookup_out;
  assign gen_inst                      = decode_inst;
  assign lookup_out                    = lut$lookup_out;
  assign lut$clk                       = clk;
  assign lut$lookup_in_[2:0]           = decode_inst[14:12];
  assign lut$reset                     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_result(rs=result_field_slice.start, re=result_field_slice.stop):
  //       s.decode_result.v = 0
  //       s.decode_result[rs:re].v = s.gen_payload

  // logic for connect_result()
  always @ (*) begin
    decode_result = 0;
    decode_result[(6)-1:0] = gen_payload;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_success():
  //       s.decode_success.v = s.gen_valid & s.and_unit.op_out

  // logic for compute_success()
  always @ (*) begin
    decode_success = (gen_valid&and_unit$op_out);
  end


endmodule // GenDecoder_0x7d917d4fc7f6270a

//-----------------------------------------------------------------------------
// LookupTable_0x3f37677ed10fc59b
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(3)) -> (valid: Bits(1), out: Bits(6))", "mapping": {"0": "func=0x0:op32=0x0:unsigned=0x0", "2": "func=0x3:op32=0x0:unsigned=0x0", "3": "func=0x3:op32=0x0:unsigned=0x1", "4": "func=0x4:op32=0x0:unsigned=0x0", "6": "func=0x7:op32=0x0:unsigned=0x0", "7": "func=0x8:op32=0x0:unsigned=0x0"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0x3f37677ed10fc59b
(
  input  logic [   0:0] clk,
  input  logic [   2:0] lookup_in_,
  output logic [   5:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   5:0] mux$mux_default;
  logic   [   5:0] mux$mux_in_$000;
  logic   [   5:0] mux$mux_in_$001;
  logic   [   5:0] mux$mux_in_$002;
  logic   [   5:0] mux$mux_in_$003;
  logic   [   5:0] mux$mux_in_$004;
  logic   [   5:0] mux$mux_in_$005;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   2:0] mux$mux_select;
  logic   [   5:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x4a721ae074151a29 mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .mux_in_$003 ( mux$mux_in_$003 ),
    .mux_in_$004 ( mux$mux_in_$004 ),
    .mux_in_$005 ( mux$mux_in_$005 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 6'd0;
  assign mux$mux_in_$000 = 6'd0;
  assign mux$mux_in_$001 = 6'd3;
  assign mux$mux_in_$002 = 6'd35;
  assign mux$mux_in_$003 = 6'd4;
  assign mux$mux_in_$004 = 6'd7;
  assign mux$mux_in_$005 = 6'd8;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0x3f37677ed10fc59b

//-----------------------------------------------------------------------------
// CaseMux_0x4a721ae074151a29
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(6), in_: Bits(6) [6], select: Bits(3)) -> (out: Bits(6), matched: Bits(1))", "svalues": ["0", "2", "3", "4", "6", "7"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x4a721ae074151a29
(
  input  logic [   0:0] clk,
  input  logic [   5:0] mux_default,
  input  logic [   5:0] mux_in_$000,
  input  logic [   5:0] mux_in_$001,
  input  logic [   5:0] mux_in_$002,
  input  logic [   5:0] mux_in_$003,
  input  logic [   5:0] mux_in_$004,
  input  logic [   5:0] mux_in_$005,
  output logic [   0:0] mux_matched,
  output logic [   5:0] mux_out,
  input  logic [   2:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   5:0] out_chain$000;
  logic   [   5:0] out_chain$001;
  logic   [   5:0] out_chain$002;
  logic   [   5:0] out_chain$003;
  logic   [   5:0] out_chain$004;
  logic   [   5:0] out_chain$005;
  logic   [   5:0] out_chain$006;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;
  logic   [   0:0] valid_chain$003;
  logic   [   0:0] valid_chain$004;
  logic   [   0:0] valid_chain$005;
  logic   [   0:0] valid_chain$006;


  // signal connections
  assign mux_matched     = valid_chain$006;
  assign mux_out         = out_chain$006;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   5:0] mux_in_[0:5];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  assign mux_in_[  3] = mux_in_$003;
  assign mux_in_[  4] = mux_in_$004;
  assign mux_in_[  5] = mux_in_$005;
  logic    [   5:0] out_chain[0:6];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  assign out_chain$003 = out_chain[  3];
  assign out_chain$004 = out_chain[  4];
  assign out_chain$005 = out_chain[  5];
  assign out_chain$006 = out_chain[  6];
  logic    [   0:0] valid_chain[0:6];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];
  assign valid_chain$003 = valid_chain[  3];
  assign valid_chain$004 = valid_chain[  4];
  assign valid_chain$005 = valid_chain[  5];
  assign valid_chain$006 = valid_chain[  6];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 0)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 2)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 3)) begin
      out_chain[3] = mux_in_[2];
      valid_chain[3] = 1;
    end
    else begin
      out_chain[3] = out_chain[2];
      valid_chain[3] = valid_chain[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 4)) begin
      out_chain[4] = mux_in_[3];
      valid_chain[4] = 1;
    end
    else begin
      out_chain[4] = out_chain[3];
      valid_chain[4] = valid_chain[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 6)) begin
      out_chain[5] = mux_in_[4];
      valid_chain[5] = 1;
    end
    else begin
      out_chain[5] = out_chain[4];
      valid_chain[5] = valid_chain[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 7)) begin
      out_chain[6] = mux_in_[5];
      valid_chain[6] = 1;
    end
    else begin
      out_chain[6] = out_chain[5];
      valid_chain[6] = valid_chain[5];
    end
  end


endmodule // CaseMux_0x4a721ae074151a29

//-----------------------------------------------------------------------------
// GenDecoderFixed_0x29e217d76d82f1af
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"ResultKind": 6, "field_list": ["funct3"], "field_map": {"0": "func=0x0:op32=0x1:unsigned=0x0"}, "fixed_map": {"opcode": "1b"}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 0, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoderFixed_0x29e217d76d82f1af
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // identity_generator temporaries
  logic   [  31:0] identity_generator$gen_inst;
  logic   [   5:0] identity_generator$gen_data;
  logic   [   0:0] identity_generator$clk;
  logic   [   0:0] identity_generator$reset;
  logic   [   5:0] identity_generator$gen_payload;
  logic   [   0:0] identity_generator$gen_valid;

  IdentityPayloadGenerator_0x6a756b13525a1482 identity_generator
  (
    .gen_inst    ( identity_generator$gen_inst ),
    .gen_data    ( identity_generator$gen_data ),
    .clk         ( identity_generator$clk ),
    .reset       ( identity_generator$reset ),
    .gen_payload ( identity_generator$gen_payload ),
    .gen_valid   ( identity_generator$gen_valid )
  );

  // decoder temporaries
  logic   [   0:0] decoder$clk;
  logic   [   5:0] decoder$gen_payload;
  logic   [  31:0] decoder$decode_inst;
  logic   [   0:0] decoder$gen_valid;
  logic   [   0:0] decoder$reset;
  logic   [  31:0] decoder$gen_inst;
  logic   [   2:0] decoder$decode_imm_type;
  logic   [   5:0] decoder$gen_data;
  logic   [   0:0] decoder$decode_serialize;
  logic   [  14:0] decoder$decode_result;
  logic   [   0:0] decoder$decode_imm_val;
  logic   [   0:0] decoder$decode_rd_val;
  logic   [   0:0] decoder$decode_rs2_val;
  logic   [   2:0] decoder$decode_op_class;
  logic   [   0:0] decoder$decode_success;
  logic   [   0:0] decoder$decode_speculative;
  logic   [   0:0] decoder$decode_rs1_val;

  GenDecoder_0x5ebc2974914a6b77 decoder
  (
    .clk                ( decoder$clk ),
    .gen_payload        ( decoder$gen_payload ),
    .decode_inst        ( decoder$decode_inst ),
    .gen_valid          ( decoder$gen_valid ),
    .reset              ( decoder$reset ),
    .gen_inst           ( decoder$gen_inst ),
    .decode_imm_type    ( decoder$decode_imm_type ),
    .gen_data           ( decoder$gen_data ),
    .decode_serialize   ( decoder$decode_serialize ),
    .decode_result      ( decoder$decode_result ),
    .decode_imm_val     ( decoder$decode_imm_val ),
    .decode_rd_val      ( decoder$decode_rd_val ),
    .decode_rs2_val     ( decoder$decode_rs2_val ),
    .decode_op_class    ( decoder$decode_op_class ),
    .decode_success     ( decoder$decode_success ),
    .decode_speculative ( decoder$decode_speculative ),
    .decode_rs1_val     ( decoder$decode_rs1_val )
  );

  // signal connections
  assign decode_imm_type             = decoder$decode_imm_type;
  assign decode_imm_val              = decoder$decode_imm_val;
  assign decode_op_class             = decoder$decode_op_class;
  assign decode_rd_val               = decoder$decode_rd_val;
  assign decode_result               = decoder$decode_result;
  assign decode_rs1_val              = decoder$decode_rs1_val;
  assign decode_rs2_val              = decoder$decode_rs2_val;
  assign decode_serialize            = decoder$decode_serialize;
  assign decode_speculative          = decoder$decode_speculative;
  assign decode_success              = decoder$decode_success;
  assign decoder$clk                 = clk;
  assign decoder$decode_inst         = decode_inst;
  assign decoder$gen_payload         = identity_generator$gen_payload;
  assign decoder$gen_valid           = identity_generator$gen_valid;
  assign decoder$reset               = reset;
  assign identity_generator$clk      = clk;
  assign identity_generator$gen_data = decoder$gen_data;
  assign identity_generator$gen_inst = decoder$gen_inst;
  assign identity_generator$reset    = reset;



endmodule // GenDecoderFixed_0x29e217d76d82f1af

//-----------------------------------------------------------------------------
// GenDecoder_0x5ebc2974914a6b77
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"In": 6, "ResultKind": 6, "field_list": ["funct3"], "field_map": {"0": "func=0x0:op32=0x1:unsigned=0x0"}, "fixed_map": {"opcode": "1b"}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 0, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoder_0x5ebc2974914a6b77
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic  [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic  [   0:0] decode_success,
  output logic [   5:0] gen_data,
  output logic [  31:0] gen_inst,
  input  logic [   5:0] gen_payload,
  input  logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] fixed_equals$000;
  logic   [   5:0] lookup_out;


  // lut temporaries
  logic   [   0:0] lut$clk;
  logic   [   0:0] lut$reset;
  logic   [   2:0] lut$lookup_in_;
  logic   [   5:0] lut$lookup_out;
  logic   [   0:0] lut$lookup_valid;

  LookupTable_0x195e36a6e48ba0db lut
  (
    .clk          ( lut$clk ),
    .reset        ( lut$reset ),
    .lookup_in_   ( lut$lookup_in_ ),
    .lookup_out   ( lut$lookup_out ),
    .lookup_valid ( lut$lookup_valid )
  );

  // equals_units$000 temporaries
  logic   [   0:0] equals_units$000$clk;
  logic   [   6:0] equals_units$000$compare_in_a;
  logic   [   6:0] equals_units$000$compare_in_b;
  logic   [   0:0] equals_units$000$reset;
  logic   [   0:0] equals_units$000$compare_out;

  Equals_0x6924ce1fe1e63d28 equals_units$000
  (
    .clk          ( equals_units$000$clk ),
    .compare_in_a ( equals_units$000$compare_in_a ),
    .compare_in_b ( equals_units$000$compare_in_b ),
    .reset        ( equals_units$000$reset ),
    .compare_out  ( equals_units$000$compare_out )
  );

  // and_unit temporaries
  logic   [   0:0] and_unit$op_in_$000;
  logic   [   0:0] and_unit$op_in_$001;
  logic   [   0:0] and_unit$clk;
  logic   [   0:0] and_unit$reset;
  logic   [   0:0] and_unit$op_out;

  And_0x8e49eae68bebab2 and_unit
  (
    .op_in_$000 ( and_unit$op_in_$000 ),
    .op_in_$001 ( and_unit$op_in_$001 ),
    .clk        ( and_unit$clk ),
    .reset      ( and_unit$reset ),
    .op_out     ( and_unit$op_out )
  );

  // signal connections
  assign and_unit$clk                  = clk;
  assign and_unit$op_in_$000           = equals_units$000$compare_out;
  assign and_unit$op_in_$001           = lut$lookup_valid;
  assign and_unit$reset                = reset;
  assign decode_imm_type               = 3'd0;
  assign decode_imm_val                = 1'd1;
  assign decode_op_class               = 3'd0;
  assign decode_rd_val                 = 1'd1;
  assign decode_rs1_val                = 1'd1;
  assign decode_rs2_val                = 1'd0;
  assign decode_serialize              = 1'd0;
  assign decode_speculative            = 1'd0;
  assign equals_units$000$clk          = clk;
  assign equals_units$000$compare_in_a = decode_inst[6:0];
  assign equals_units$000$compare_in_b = 7'd27;
  assign equals_units$000$reset        = reset;
  assign gen_data                      = lookup_out;
  assign gen_inst                      = decode_inst;
  assign lookup_out                    = lut$lookup_out;
  assign lut$clk                       = clk;
  assign lut$lookup_in_[2:0]           = decode_inst[14:12];
  assign lut$reset                     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_result(rs=result_field_slice.start, re=result_field_slice.stop):
  //       s.decode_result.v = 0
  //       s.decode_result[rs:re].v = s.gen_payload

  // logic for connect_result()
  always @ (*) begin
    decode_result = 0;
    decode_result[(6)-1:0] = gen_payload;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_success():
  //       s.decode_success.v = s.gen_valid & s.and_unit.op_out

  // logic for compute_success()
  always @ (*) begin
    decode_success = (gen_valid&and_unit$op_out);
  end


endmodule // GenDecoder_0x5ebc2974914a6b77

//-----------------------------------------------------------------------------
// LookupTable_0x195e36a6e48ba0db
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(3)) -> (valid: Bits(1), out: Bits(6))", "mapping": {"0": "func=0x0:op32=0x1:unsigned=0x0"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0x195e36a6e48ba0db
(
  input  logic [   0:0] clk,
  input  logic [   2:0] lookup_in_,
  output logic [   5:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   5:0] mux$mux_default;
  logic   [   5:0] mux$mux_in_$000;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   2:0] mux$mux_select;
  logic   [   5:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x325c3116b59e5559 mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 6'd0;
  assign mux$mux_in_$000 = 6'd16;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0x195e36a6e48ba0db

//-----------------------------------------------------------------------------
// CaseMux_0x325c3116b59e5559
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(6), in_: Bits(6) [1], select: Bits(3)) -> (out: Bits(6), matched: Bits(1))", "svalues": ["0"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x325c3116b59e5559
(
  input  logic [   0:0] clk,
  input  logic [   5:0] mux_default,
  input  logic [   5:0] mux_in_$000,
  output logic [   0:0] mux_matched,
  output logic [   5:0] mux_out,
  input  logic [   2:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   5:0] out_chain$000;
  logic   [   5:0] out_chain$001;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;


  // signal connections
  assign mux_matched     = valid_chain$001;
  assign mux_out         = out_chain$001;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   5:0] mux_in_[0:0];
  assign mux_in_[  0] = mux_in_$000;
  logic    [   5:0] out_chain[0:1];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  logic    [   0:0] valid_chain[0:1];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 0)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end


endmodule // CaseMux_0x325c3116b59e5559

//-----------------------------------------------------------------------------
// GenDecoderFixed_0x2f940af682bd257
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"ResultKind": 6, "field_list": ["funct7_shft64", "funct3"], "field_map": {"(0, 1)": "func=0x2:op32=0x0:unsigned=0x0", "(0, 5)": "func=0x5:op32=0x0:unsigned=0x0", "(16, 5)": "func=0x6:op32=0x0:unsigned=0x0"}, "fixed_map": {"opcode": "13"}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 0, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoderFixed_0x2f940af682bd257
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // identity_generator temporaries
  logic   [  31:0] identity_generator$gen_inst;
  logic   [   5:0] identity_generator$gen_data;
  logic   [   0:0] identity_generator$clk;
  logic   [   0:0] identity_generator$reset;
  logic   [   5:0] identity_generator$gen_payload;
  logic   [   0:0] identity_generator$gen_valid;

  IdentityPayloadGenerator_0x6a756b13525a1482 identity_generator
  (
    .gen_inst    ( identity_generator$gen_inst ),
    .gen_data    ( identity_generator$gen_data ),
    .clk         ( identity_generator$clk ),
    .reset       ( identity_generator$reset ),
    .gen_payload ( identity_generator$gen_payload ),
    .gen_valid   ( identity_generator$gen_valid )
  );

  // decoder temporaries
  logic   [   0:0] decoder$clk;
  logic   [   5:0] decoder$gen_payload;
  logic   [  31:0] decoder$decode_inst;
  logic   [   0:0] decoder$gen_valid;
  logic   [   0:0] decoder$reset;
  logic   [  31:0] decoder$gen_inst;
  logic   [   2:0] decoder$decode_imm_type;
  logic   [   5:0] decoder$gen_data;
  logic   [   0:0] decoder$decode_serialize;
  logic   [  14:0] decoder$decode_result;
  logic   [   0:0] decoder$decode_imm_val;
  logic   [   0:0] decoder$decode_rd_val;
  logic   [   0:0] decoder$decode_rs2_val;
  logic   [   2:0] decoder$decode_op_class;
  logic   [   0:0] decoder$decode_success;
  logic   [   0:0] decoder$decode_speculative;
  logic   [   0:0] decoder$decode_rs1_val;

  GenDecoder_0x3c9b01c59fa9386b decoder
  (
    .clk                ( decoder$clk ),
    .gen_payload        ( decoder$gen_payload ),
    .decode_inst        ( decoder$decode_inst ),
    .gen_valid          ( decoder$gen_valid ),
    .reset              ( decoder$reset ),
    .gen_inst           ( decoder$gen_inst ),
    .decode_imm_type    ( decoder$decode_imm_type ),
    .gen_data           ( decoder$gen_data ),
    .decode_serialize   ( decoder$decode_serialize ),
    .decode_result      ( decoder$decode_result ),
    .decode_imm_val     ( decoder$decode_imm_val ),
    .decode_rd_val      ( decoder$decode_rd_val ),
    .decode_rs2_val     ( decoder$decode_rs2_val ),
    .decode_op_class    ( decoder$decode_op_class ),
    .decode_success     ( decoder$decode_success ),
    .decode_speculative ( decoder$decode_speculative ),
    .decode_rs1_val     ( decoder$decode_rs1_val )
  );

  // signal connections
  assign decode_imm_type             = decoder$decode_imm_type;
  assign decode_imm_val              = decoder$decode_imm_val;
  assign decode_op_class             = decoder$decode_op_class;
  assign decode_rd_val               = decoder$decode_rd_val;
  assign decode_result               = decoder$decode_result;
  assign decode_rs1_val              = decoder$decode_rs1_val;
  assign decode_rs2_val              = decoder$decode_rs2_val;
  assign decode_serialize            = decoder$decode_serialize;
  assign decode_speculative          = decoder$decode_speculative;
  assign decode_success              = decoder$decode_success;
  assign decoder$clk                 = clk;
  assign decoder$decode_inst         = decode_inst;
  assign decoder$gen_payload         = identity_generator$gen_payload;
  assign decoder$gen_valid           = identity_generator$gen_valid;
  assign decoder$reset               = reset;
  assign identity_generator$clk      = clk;
  assign identity_generator$gen_data = decoder$gen_data;
  assign identity_generator$gen_inst = decoder$gen_inst;
  assign identity_generator$reset    = reset;



endmodule // GenDecoderFixed_0x2f940af682bd257

//-----------------------------------------------------------------------------
// GenDecoder_0x3c9b01c59fa9386b
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"In": 6, "ResultKind": 6, "field_list": ["funct7_shft64", "funct3"], "field_map": {"(0, 1)": "func=0x2:op32=0x0:unsigned=0x0", "(0, 5)": "func=0x5:op32=0x0:unsigned=0x0", "(16, 5)": "func=0x6:op32=0x0:unsigned=0x0"}, "fixed_map": {"opcode": "13"}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 0, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoder_0x3c9b01c59fa9386b
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic  [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic  [   0:0] decode_success,
  output logic [   5:0] gen_data,
  output logic [  31:0] gen_inst,
  input  logic [   5:0] gen_payload,
  input  logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] fixed_equals$000;
  logic   [   5:0] lookup_out;


  // lut temporaries
  logic   [   0:0] lut$clk;
  logic   [   0:0] lut$reset;
  logic   [   8:0] lut$lookup_in_;
  logic   [   5:0] lut$lookup_out;
  logic   [   0:0] lut$lookup_valid;

  LookupTable_0x577585e517feb282 lut
  (
    .clk          ( lut$clk ),
    .reset        ( lut$reset ),
    .lookup_in_   ( lut$lookup_in_ ),
    .lookup_out   ( lut$lookup_out ),
    .lookup_valid ( lut$lookup_valid )
  );

  // equals_units$000 temporaries
  logic   [   0:0] equals_units$000$clk;
  logic   [   6:0] equals_units$000$compare_in_a;
  logic   [   6:0] equals_units$000$compare_in_b;
  logic   [   0:0] equals_units$000$reset;
  logic   [   0:0] equals_units$000$compare_out;

  Equals_0x6924ce1fe1e63d28 equals_units$000
  (
    .clk          ( equals_units$000$clk ),
    .compare_in_a ( equals_units$000$compare_in_a ),
    .compare_in_b ( equals_units$000$compare_in_b ),
    .reset        ( equals_units$000$reset ),
    .compare_out  ( equals_units$000$compare_out )
  );

  // and_unit temporaries
  logic   [   0:0] and_unit$op_in_$000;
  logic   [   0:0] and_unit$op_in_$001;
  logic   [   0:0] and_unit$clk;
  logic   [   0:0] and_unit$reset;
  logic   [   0:0] and_unit$op_out;

  And_0x8e49eae68bebab2 and_unit
  (
    .op_in_$000 ( and_unit$op_in_$000 ),
    .op_in_$001 ( and_unit$op_in_$001 ),
    .clk        ( and_unit$clk ),
    .reset      ( and_unit$reset ),
    .op_out     ( and_unit$op_out )
  );

  // signal connections
  assign and_unit$clk                  = clk;
  assign and_unit$op_in_$000           = equals_units$000$compare_out;
  assign and_unit$op_in_$001           = lut$lookup_valid;
  assign and_unit$reset                = reset;
  assign decode_imm_type               = 3'd7;
  assign decode_imm_val                = 1'd1;
  assign decode_op_class               = 3'd0;
  assign decode_rd_val                 = 1'd1;
  assign decode_rs1_val                = 1'd1;
  assign decode_rs2_val                = 1'd0;
  assign decode_serialize              = 1'd0;
  assign decode_speculative            = 1'd0;
  assign equals_units$000$clk          = clk;
  assign equals_units$000$compare_in_a = decode_inst[6:0];
  assign equals_units$000$compare_in_b = 7'd19;
  assign equals_units$000$reset        = reset;
  assign gen_data                      = lookup_out;
  assign gen_inst                      = decode_inst;
  assign lookup_out                    = lut$lookup_out;
  assign lut$clk                       = clk;
  assign lut$lookup_in_[5:0]           = decode_inst[31:26];
  assign lut$lookup_in_[8:6]           = decode_inst[14:12];
  assign lut$reset                     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_result(rs=result_field_slice.start, re=result_field_slice.stop):
  //       s.decode_result.v = 0
  //       s.decode_result[rs:re].v = s.gen_payload

  // logic for connect_result()
  always @ (*) begin
    decode_result = 0;
    decode_result[(6)-1:0] = gen_payload;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_success():
  //       s.decode_success.v = s.gen_valid & s.and_unit.op_out

  // logic for compute_success()
  always @ (*) begin
    decode_success = (gen_valid&and_unit$op_out);
  end


endmodule // GenDecoder_0x3c9b01c59fa9386b

//-----------------------------------------------------------------------------
// LookupTable_0x577585e517feb282
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(9)) -> (valid: Bits(1), out: Bits(6))", "mapping": {"040": "func=0x2:op32=0x0:unsigned=0x0", "140": "func=0x5:op32=0x0:unsigned=0x0", "150": "func=0x6:op32=0x0:unsigned=0x0"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0x577585e517feb282
(
  input  logic [   0:0] clk,
  input  logic [   8:0] lookup_in_,
  output logic [   5:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   5:0] mux$mux_default;
  logic   [   5:0] mux$mux_in_$000;
  logic   [   5:0] mux$mux_in_$001;
  logic   [   5:0] mux$mux_in_$002;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   8:0] mux$mux_select;
  logic   [   5:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x5acffc90b50b40c0 mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 6'd0;
  assign mux$mux_in_$000 = 6'd2;
  assign mux$mux_in_$001 = 6'd5;
  assign mux$mux_in_$002 = 6'd6;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0x577585e517feb282

//-----------------------------------------------------------------------------
// CaseMux_0x5acffc90b50b40c0
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(6), in_: Bits(6) [3], select: Bits(9)) -> (out: Bits(6), matched: Bits(1))", "svalues": ["040", "140", "150"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x5acffc90b50b40c0
(
  input  logic [   0:0] clk,
  input  logic [   5:0] mux_default,
  input  logic [   5:0] mux_in_$000,
  input  logic [   5:0] mux_in_$001,
  input  logic [   5:0] mux_in_$002,
  output logic [   0:0] mux_matched,
  output logic [   5:0] mux_out,
  input  logic [   8:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   5:0] out_chain$000;
  logic   [   5:0] out_chain$001;
  logic   [   5:0] out_chain$002;
  logic   [   5:0] out_chain$003;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;
  logic   [   0:0] valid_chain$003;


  // signal connections
  assign mux_matched     = valid_chain$003;
  assign mux_out         = out_chain$003;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   5:0] mux_in_[0:2];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  logic    [   5:0] out_chain[0:3];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  assign out_chain$003 = out_chain[  3];
  logic    [   0:0] valid_chain[0:3];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];
  assign valid_chain$003 = valid_chain[  3];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 64)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 320)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 336)) begin
      out_chain[3] = mux_in_[2];
      valid_chain[3] = 1;
    end
    else begin
      out_chain[3] = out_chain[2];
      valid_chain[3] = valid_chain[2];
    end
  end


endmodule // CaseMux_0x5acffc90b50b40c0

//-----------------------------------------------------------------------------
// GenDecoderFixed_0x55d6eb7561f62d2e
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"ResultKind": 6, "field_list": ["funct7", "funct3"], "field_map": {"(0, 1)": "func=0x2:op32=0x1:unsigned=0x0", "(0, 5)": "func=0x5:op32=0x1:unsigned=0x0", "(32, 5)": "func=0x6:op32=0x1:unsigned=0x0"}, "fixed_map": {"opcode": "1b"}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 0, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoderFixed_0x55d6eb7561f62d2e
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // identity_generator temporaries
  logic   [  31:0] identity_generator$gen_inst;
  logic   [   5:0] identity_generator$gen_data;
  logic   [   0:0] identity_generator$clk;
  logic   [   0:0] identity_generator$reset;
  logic   [   5:0] identity_generator$gen_payload;
  logic   [   0:0] identity_generator$gen_valid;

  IdentityPayloadGenerator_0x6a756b13525a1482 identity_generator
  (
    .gen_inst    ( identity_generator$gen_inst ),
    .gen_data    ( identity_generator$gen_data ),
    .clk         ( identity_generator$clk ),
    .reset       ( identity_generator$reset ),
    .gen_payload ( identity_generator$gen_payload ),
    .gen_valid   ( identity_generator$gen_valid )
  );

  // decoder temporaries
  logic   [   0:0] decoder$clk;
  logic   [   5:0] decoder$gen_payload;
  logic   [  31:0] decoder$decode_inst;
  logic   [   0:0] decoder$gen_valid;
  logic   [   0:0] decoder$reset;
  logic   [  31:0] decoder$gen_inst;
  logic   [   2:0] decoder$decode_imm_type;
  logic   [   5:0] decoder$gen_data;
  logic   [   0:0] decoder$decode_serialize;
  logic   [  14:0] decoder$decode_result;
  logic   [   0:0] decoder$decode_imm_val;
  logic   [   0:0] decoder$decode_rd_val;
  logic   [   0:0] decoder$decode_rs2_val;
  logic   [   2:0] decoder$decode_op_class;
  logic   [   0:0] decoder$decode_success;
  logic   [   0:0] decoder$decode_speculative;
  logic   [   0:0] decoder$decode_rs1_val;

  GenDecoder_0x67895dbf831f0886 decoder
  (
    .clk                ( decoder$clk ),
    .gen_payload        ( decoder$gen_payload ),
    .decode_inst        ( decoder$decode_inst ),
    .gen_valid          ( decoder$gen_valid ),
    .reset              ( decoder$reset ),
    .gen_inst           ( decoder$gen_inst ),
    .decode_imm_type    ( decoder$decode_imm_type ),
    .gen_data           ( decoder$gen_data ),
    .decode_serialize   ( decoder$decode_serialize ),
    .decode_result      ( decoder$decode_result ),
    .decode_imm_val     ( decoder$decode_imm_val ),
    .decode_rd_val      ( decoder$decode_rd_val ),
    .decode_rs2_val     ( decoder$decode_rs2_val ),
    .decode_op_class    ( decoder$decode_op_class ),
    .decode_success     ( decoder$decode_success ),
    .decode_speculative ( decoder$decode_speculative ),
    .decode_rs1_val     ( decoder$decode_rs1_val )
  );

  // signal connections
  assign decode_imm_type             = decoder$decode_imm_type;
  assign decode_imm_val              = decoder$decode_imm_val;
  assign decode_op_class             = decoder$decode_op_class;
  assign decode_rd_val               = decoder$decode_rd_val;
  assign decode_result               = decoder$decode_result;
  assign decode_rs1_val              = decoder$decode_rs1_val;
  assign decode_rs2_val              = decoder$decode_rs2_val;
  assign decode_serialize            = decoder$decode_serialize;
  assign decode_speculative          = decoder$decode_speculative;
  assign decode_success              = decoder$decode_success;
  assign decoder$clk                 = clk;
  assign decoder$decode_inst         = decode_inst;
  assign decoder$gen_payload         = identity_generator$gen_payload;
  assign decoder$gen_valid           = identity_generator$gen_valid;
  assign decoder$reset               = reset;
  assign identity_generator$clk      = clk;
  assign identity_generator$gen_data = decoder$gen_data;
  assign identity_generator$gen_inst = decoder$gen_inst;
  assign identity_generator$reset    = reset;



endmodule // GenDecoderFixed_0x55d6eb7561f62d2e

//-----------------------------------------------------------------------------
// GenDecoder_0x67895dbf831f0886
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"In": 6, "ResultKind": 6, "field_list": ["funct7", "funct3"], "field_map": {"(0, 1)": "func=0x2:op32=0x1:unsigned=0x0", "(0, 5)": "func=0x5:op32=0x1:unsigned=0x0", "(32, 5)": "func=0x6:op32=0x1:unsigned=0x0"}, "fixed_map": {"opcode": "1b"}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 1, "rs2_val": 0, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoder_0x67895dbf831f0886
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic  [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic  [   0:0] decode_success,
  output logic [   5:0] gen_data,
  output logic [  31:0] gen_inst,
  input  logic [   5:0] gen_payload,
  input  logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] fixed_equals$000;
  logic   [   5:0] lookup_out;


  // lut temporaries
  logic   [   0:0] lut$clk;
  logic   [   0:0] lut$reset;
  logic   [   9:0] lut$lookup_in_;
  logic   [   5:0] lut$lookup_out;
  logic   [   0:0] lut$lookup_valid;

  LookupTable_0x72ea311964667966 lut
  (
    .clk          ( lut$clk ),
    .reset        ( lut$reset ),
    .lookup_in_   ( lut$lookup_in_ ),
    .lookup_out   ( lut$lookup_out ),
    .lookup_valid ( lut$lookup_valid )
  );

  // equals_units$000 temporaries
  logic   [   0:0] equals_units$000$clk;
  logic   [   6:0] equals_units$000$compare_in_a;
  logic   [   6:0] equals_units$000$compare_in_b;
  logic   [   0:0] equals_units$000$reset;
  logic   [   0:0] equals_units$000$compare_out;

  Equals_0x6924ce1fe1e63d28 equals_units$000
  (
    .clk          ( equals_units$000$clk ),
    .compare_in_a ( equals_units$000$compare_in_a ),
    .compare_in_b ( equals_units$000$compare_in_b ),
    .reset        ( equals_units$000$reset ),
    .compare_out  ( equals_units$000$compare_out )
  );

  // and_unit temporaries
  logic   [   0:0] and_unit$op_in_$000;
  logic   [   0:0] and_unit$op_in_$001;
  logic   [   0:0] and_unit$clk;
  logic   [   0:0] and_unit$reset;
  logic   [   0:0] and_unit$op_out;

  And_0x8e49eae68bebab2 and_unit
  (
    .op_in_$000 ( and_unit$op_in_$000 ),
    .op_in_$001 ( and_unit$op_in_$001 ),
    .clk        ( and_unit$clk ),
    .reset      ( and_unit$reset ),
    .op_out     ( and_unit$op_out )
  );

  // signal connections
  assign and_unit$clk                  = clk;
  assign and_unit$op_in_$000           = equals_units$000$compare_out;
  assign and_unit$op_in_$001           = lut$lookup_valid;
  assign and_unit$reset                = reset;
  assign decode_imm_type               = 3'd7;
  assign decode_imm_val                = 1'd1;
  assign decode_op_class               = 3'd0;
  assign decode_rd_val                 = 1'd1;
  assign decode_rs1_val                = 1'd1;
  assign decode_rs2_val                = 1'd0;
  assign decode_serialize              = 1'd0;
  assign decode_speculative            = 1'd0;
  assign equals_units$000$clk          = clk;
  assign equals_units$000$compare_in_a = decode_inst[6:0];
  assign equals_units$000$compare_in_b = 7'd27;
  assign equals_units$000$reset        = reset;
  assign gen_data                      = lookup_out;
  assign gen_inst                      = decode_inst;
  assign lookup_out                    = lut$lookup_out;
  assign lut$clk                       = clk;
  assign lut$lookup_in_[6:0]           = decode_inst[31:25];
  assign lut$lookup_in_[9:7]           = decode_inst[14:12];
  assign lut$reset                     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_result(rs=result_field_slice.start, re=result_field_slice.stop):
  //       s.decode_result.v = 0
  //       s.decode_result[rs:re].v = s.gen_payload

  // logic for connect_result()
  always @ (*) begin
    decode_result = 0;
    decode_result[(6)-1:0] = gen_payload;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_success():
  //       s.decode_success.v = s.gen_valid & s.and_unit.op_out

  // logic for compute_success()
  always @ (*) begin
    decode_success = (gen_valid&and_unit$op_out);
  end


endmodule // GenDecoder_0x67895dbf831f0886

//-----------------------------------------------------------------------------
// LookupTable_0x72ea311964667966
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(10)) -> (valid: Bits(1), out: Bits(6))", "mapping": {"080": "func=0x2:op32=0x1:unsigned=0x0", "280": "func=0x5:op32=0x1:unsigned=0x0", "2a0": "func=0x6:op32=0x1:unsigned=0x0"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0x72ea311964667966
(
  input  logic [   0:0] clk,
  input  logic [   9:0] lookup_in_,
  output logic [   5:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   5:0] mux$mux_default;
  logic   [   5:0] mux$mux_in_$000;
  logic   [   5:0] mux$mux_in_$001;
  logic   [   5:0] mux$mux_in_$002;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   9:0] mux$mux_select;
  logic   [   5:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x42488f7e692de783 mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 6'd0;
  assign mux$mux_in_$000 = 6'd18;
  assign mux$mux_in_$001 = 6'd21;
  assign mux$mux_in_$002 = 6'd22;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0x72ea311964667966

//-----------------------------------------------------------------------------
// CaseMux_0x42488f7e692de783
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(6), in_: Bits(6) [3], select: Bits(10)) -> (out: Bits(6), matched: Bits(1))", "svalues": ["080", "280", "2a0"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x42488f7e692de783
(
  input  logic [   0:0] clk,
  input  logic [   5:0] mux_default,
  input  logic [   5:0] mux_in_$000,
  input  logic [   5:0] mux_in_$001,
  input  logic [   5:0] mux_in_$002,
  output logic [   0:0] mux_matched,
  output logic [   5:0] mux_out,
  input  logic [   9:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   5:0] out_chain$000;
  logic   [   5:0] out_chain$001;
  logic   [   5:0] out_chain$002;
  logic   [   5:0] out_chain$003;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;
  logic   [   0:0] valid_chain$003;


  // signal connections
  assign mux_matched     = valid_chain$003;
  assign mux_out         = out_chain$003;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   5:0] mux_in_[0:2];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  logic    [   5:0] out_chain[0:3];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  assign out_chain$003 = out_chain[  3];
  logic    [   0:0] valid_chain[0:3];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];
  assign valid_chain$003 = valid_chain[  3];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 128)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 640)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 672)) begin
      out_chain[3] = mux_in_[2];
      valid_chain[3] = 1;
    end
    else begin
      out_chain[3] = out_chain[2];
      valid_chain[3] = valid_chain[2];
    end
  end


endmodule // CaseMux_0x42488f7e692de783

//-----------------------------------------------------------------------------
// GenDecoderFixed_0x33541dea129c9660
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"ResultKind": 6, "field_list": ["opcode"], "field_map": {"17": "func=0xa:op32=0x0:unsigned=0x0", "37": "func=0x9:op32=0x0:unsigned=0x0"}, "fixed_map": {}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 0, "rs2_val": 0, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoderFixed_0x33541dea129c9660
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // identity_generator temporaries
  logic   [  31:0] identity_generator$gen_inst;
  logic   [   5:0] identity_generator$gen_data;
  logic   [   0:0] identity_generator$clk;
  logic   [   0:0] identity_generator$reset;
  logic   [   5:0] identity_generator$gen_payload;
  logic   [   0:0] identity_generator$gen_valid;

  IdentityPayloadGenerator_0x6a756b13525a1482 identity_generator
  (
    .gen_inst    ( identity_generator$gen_inst ),
    .gen_data    ( identity_generator$gen_data ),
    .clk         ( identity_generator$clk ),
    .reset       ( identity_generator$reset ),
    .gen_payload ( identity_generator$gen_payload ),
    .gen_valid   ( identity_generator$gen_valid )
  );

  // decoder temporaries
  logic   [   0:0] decoder$clk;
  logic   [   5:0] decoder$gen_payload;
  logic   [  31:0] decoder$decode_inst;
  logic   [   0:0] decoder$gen_valid;
  logic   [   0:0] decoder$reset;
  logic   [  31:0] decoder$gen_inst;
  logic   [   2:0] decoder$decode_imm_type;
  logic   [   5:0] decoder$gen_data;
  logic   [   0:0] decoder$decode_serialize;
  logic   [  14:0] decoder$decode_result;
  logic   [   0:0] decoder$decode_imm_val;
  logic   [   0:0] decoder$decode_rd_val;
  logic   [   0:0] decoder$decode_rs2_val;
  logic   [   2:0] decoder$decode_op_class;
  logic   [   0:0] decoder$decode_success;
  logic   [   0:0] decoder$decode_speculative;
  logic   [   0:0] decoder$decode_rs1_val;

  GenDecoder_0x5eeb8a1ab37ed9c4 decoder
  (
    .clk                ( decoder$clk ),
    .gen_payload        ( decoder$gen_payload ),
    .decode_inst        ( decoder$decode_inst ),
    .gen_valid          ( decoder$gen_valid ),
    .reset              ( decoder$reset ),
    .gen_inst           ( decoder$gen_inst ),
    .decode_imm_type    ( decoder$decode_imm_type ),
    .gen_data           ( decoder$gen_data ),
    .decode_serialize   ( decoder$decode_serialize ),
    .decode_result      ( decoder$decode_result ),
    .decode_imm_val     ( decoder$decode_imm_val ),
    .decode_rd_val      ( decoder$decode_rd_val ),
    .decode_rs2_val     ( decoder$decode_rs2_val ),
    .decode_op_class    ( decoder$decode_op_class ),
    .decode_success     ( decoder$decode_success ),
    .decode_speculative ( decoder$decode_speculative ),
    .decode_rs1_val     ( decoder$decode_rs1_val )
  );

  // signal connections
  assign decode_imm_type             = decoder$decode_imm_type;
  assign decode_imm_val              = decoder$decode_imm_val;
  assign decode_op_class             = decoder$decode_op_class;
  assign decode_rd_val               = decoder$decode_rd_val;
  assign decode_result               = decoder$decode_result;
  assign decode_rs1_val              = decoder$decode_rs1_val;
  assign decode_rs2_val              = decoder$decode_rs2_val;
  assign decode_serialize            = decoder$decode_serialize;
  assign decode_speculative          = decoder$decode_speculative;
  assign decode_success              = decoder$decode_success;
  assign decoder$clk                 = clk;
  assign decoder$decode_inst         = decode_inst;
  assign decoder$gen_payload         = identity_generator$gen_payload;
  assign decoder$gen_valid           = identity_generator$gen_valid;
  assign decoder$reset               = reset;
  assign identity_generator$clk      = clk;
  assign identity_generator$gen_data = decoder$gen_data;
  assign identity_generator$gen_inst = decoder$gen_inst;
  assign identity_generator$reset    = reset;



endmodule // GenDecoderFixed_0x33541dea129c9660

//-----------------------------------------------------------------------------
// GenDecoder_0x5eeb8a1ab37ed9c4
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"In": 6, "ResultKind": 6, "field_list": ["opcode"], "field_map": {"17": "func=0xa:op32=0x0:unsigned=0x0", "37": "func=0x9:op32=0x0:unsigned=0x0"}, "fixed_map": {}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 1, "result_field": "alu_msg", "rs1_val": 0, "rs2_val": 0, "serialize": 0, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoder_0x5eeb8a1ab37ed9c4
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic  [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic  [   0:0] decode_success,
  output logic [   5:0] gen_data,
  output logic [  31:0] gen_inst,
  input  logic [   5:0] gen_payload,
  input  logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   5:0] lookup_out;


  // lut temporaries
  logic   [   0:0] lut$clk;
  logic   [   0:0] lut$reset;
  logic   [   6:0] lut$lookup_in_;
  logic   [   5:0] lut$lookup_out;
  logic   [   0:0] lut$lookup_valid;

  LookupTable_0x7c2fc2f3fed0bf31 lut
  (
    .clk          ( lut$clk ),
    .reset        ( lut$reset ),
    .lookup_in_   ( lut$lookup_in_ ),
    .lookup_out   ( lut$lookup_out ),
    .lookup_valid ( lut$lookup_valid )
  );

  // and_unit temporaries
  logic   [   0:0] and_unit$op_in_$000;
  logic   [   0:0] and_unit$clk;
  logic   [   0:0] and_unit$reset;
  logic   [   0:0] and_unit$op_out;

  And_0x470fbdee6c6763c5 and_unit
  (
    .op_in_$000 ( and_unit$op_in_$000 ),
    .clk        ( and_unit$clk ),
    .reset      ( and_unit$reset ),
    .op_out     ( and_unit$op_out )
  );

  // signal connections
  assign and_unit$clk        = clk;
  assign and_unit$op_in_$000 = lut$lookup_valid;
  assign and_unit$reset      = reset;
  assign decode_imm_type     = 3'd3;
  assign decode_imm_val      = 1'd1;
  assign decode_op_class     = 3'd0;
  assign decode_rd_val       = 1'd1;
  assign decode_rs1_val      = 1'd0;
  assign decode_rs2_val      = 1'd0;
  assign decode_serialize    = 1'd0;
  assign decode_speculative  = 1'd0;
  assign gen_data            = lookup_out;
  assign gen_inst            = decode_inst;
  assign lookup_out          = lut$lookup_out;
  assign lut$clk             = clk;
  assign lut$lookup_in_[6:0] = decode_inst[6:0];
  assign lut$reset           = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_result(rs=result_field_slice.start, re=result_field_slice.stop):
  //       s.decode_result.v = 0
  //       s.decode_result[rs:re].v = s.gen_payload

  // logic for connect_result()
  always @ (*) begin
    decode_result = 0;
    decode_result[(6)-1:0] = gen_payload;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_success():
  //       s.decode_success.v = s.gen_valid & s.and_unit.op_out

  // logic for compute_success()
  always @ (*) begin
    decode_success = (gen_valid&and_unit$op_out);
  end


endmodule // GenDecoder_0x5eeb8a1ab37ed9c4

//-----------------------------------------------------------------------------
// LookupTable_0x7c2fc2f3fed0bf31
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(7)) -> (valid: Bits(1), out: Bits(6))", "mapping": {"17": "func=0xa:op32=0x0:unsigned=0x0", "37": "func=0x9:op32=0x0:unsigned=0x0"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0x7c2fc2f3fed0bf31
(
  input  logic [   0:0] clk,
  input  logic [   6:0] lookup_in_,
  output logic [   5:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   5:0] mux$mux_default;
  logic   [   5:0] mux$mux_in_$000;
  logic   [   5:0] mux$mux_in_$001;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   6:0] mux$mux_select;
  logic   [   5:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x6c3b0e8f937dcf59 mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 6'd0;
  assign mux$mux_in_$000 = 6'd10;
  assign mux$mux_in_$001 = 6'd9;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0x7c2fc2f3fed0bf31

//-----------------------------------------------------------------------------
// CaseMux_0x6c3b0e8f937dcf59
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(6), in_: Bits(6) [2], select: Bits(7)) -> (out: Bits(6), matched: Bits(1))", "svalues": ["17", "37"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x6c3b0e8f937dcf59
(
  input  logic [   0:0] clk,
  input  logic [   5:0] mux_default,
  input  logic [   5:0] mux_in_$000,
  input  logic [   5:0] mux_in_$001,
  output logic [   0:0] mux_matched,
  output logic [   5:0] mux_out,
  input  logic [   6:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   5:0] out_chain$000;
  logic   [   5:0] out_chain$001;
  logic   [   5:0] out_chain$002;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;


  // signal connections
  assign mux_matched     = valid_chain$002;
  assign mux_out         = out_chain$002;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   5:0] mux_in_[0:1];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  logic    [   5:0] out_chain[0:2];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  logic    [   0:0] valid_chain[0:2];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 23)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 55)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end


endmodule // CaseMux_0x6c3b0e8f937dcf59

//-----------------------------------------------------------------------------
// And_0x470fbdee6c6763c5
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.logic {"interface": "op (in_: Bits(1) [1]) -> (out: Bits(1))"}
// PyMTL: verilator_xinit = zeros
module And_0x470fbdee6c6763c5
(
  input  logic [   0:0] clk,
  input  logic [   0:0] op_in_$000,
  output logic [   0:0] op_out,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] partials$000;


  // signal connections
  assign op_out = partials$000;

  // array declarations
  logic   [   0:0] op_in_[0:0];
  assign op_in_[  0] = op_in_$000;
  logic    [   0:0] partials[0:0];
  assign partials$000 = partials[  0];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def initial():
  //           s.partials[0].v = s.op_in_[0]

  // logic for initial()
  always @ (*) begin
    partials[0] = op_in_[0];
  end


endmodule // And_0x470fbdee6c6763c5

//-----------------------------------------------------------------------------
// CompositeDecoder_0x2c27817f254c2cc0
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"nchildren": 7}
// PyMTL: verilator_xinit = zeros
module CompositeDecoder_0x2c27817f254c2cc0
(
  input  logic [   0:0] clk,
  input  logic [   2:0] decode_child_imm_type$000,
  input  logic [   2:0] decode_child_imm_type$001,
  input  logic [   2:0] decode_child_imm_type$002,
  input  logic [   2:0] decode_child_imm_type$003,
  input  logic [   2:0] decode_child_imm_type$004,
  input  logic [   2:0] decode_child_imm_type$005,
  input  logic [   2:0] decode_child_imm_type$006,
  input  logic [   0:0] decode_child_imm_val$000,
  input  logic [   0:0] decode_child_imm_val$001,
  input  logic [   0:0] decode_child_imm_val$002,
  input  logic [   0:0] decode_child_imm_val$003,
  input  logic [   0:0] decode_child_imm_val$004,
  input  logic [   0:0] decode_child_imm_val$005,
  input  logic [   0:0] decode_child_imm_val$006,
  output logic [  31:0] decode_child_inst$000,
  output logic [  31:0] decode_child_inst$001,
  output logic [  31:0] decode_child_inst$002,
  output logic [  31:0] decode_child_inst$003,
  output logic [  31:0] decode_child_inst$004,
  output logic [  31:0] decode_child_inst$005,
  output logic [  31:0] decode_child_inst$006,
  input  logic [   2:0] decode_child_op_class$000,
  input  logic [   2:0] decode_child_op_class$001,
  input  logic [   2:0] decode_child_op_class$002,
  input  logic [   2:0] decode_child_op_class$003,
  input  logic [   2:0] decode_child_op_class$004,
  input  logic [   2:0] decode_child_op_class$005,
  input  logic [   2:0] decode_child_op_class$006,
  input  logic [   0:0] decode_child_rd_val$000,
  input  logic [   0:0] decode_child_rd_val$001,
  input  logic [   0:0] decode_child_rd_val$002,
  input  logic [   0:0] decode_child_rd_val$003,
  input  logic [   0:0] decode_child_rd_val$004,
  input  logic [   0:0] decode_child_rd_val$005,
  input  logic [   0:0] decode_child_rd_val$006,
  input  logic [  14:0] decode_child_result$000,
  input  logic [  14:0] decode_child_result$001,
  input  logic [  14:0] decode_child_result$002,
  input  logic [  14:0] decode_child_result$003,
  input  logic [  14:0] decode_child_result$004,
  input  logic [  14:0] decode_child_result$005,
  input  logic [  14:0] decode_child_result$006,
  input  logic [   0:0] decode_child_rs1_val$000,
  input  logic [   0:0] decode_child_rs1_val$001,
  input  logic [   0:0] decode_child_rs1_val$002,
  input  logic [   0:0] decode_child_rs1_val$003,
  input  logic [   0:0] decode_child_rs1_val$004,
  input  logic [   0:0] decode_child_rs1_val$005,
  input  logic [   0:0] decode_child_rs1_val$006,
  input  logic [   0:0] decode_child_rs2_val$000,
  input  logic [   0:0] decode_child_rs2_val$001,
  input  logic [   0:0] decode_child_rs2_val$002,
  input  logic [   0:0] decode_child_rs2_val$003,
  input  logic [   0:0] decode_child_rs2_val$004,
  input  logic [   0:0] decode_child_rs2_val$005,
  input  logic [   0:0] decode_child_rs2_val$006,
  input  logic [   0:0] decode_child_serialize$000,
  input  logic [   0:0] decode_child_serialize$001,
  input  logic [   0:0] decode_child_serialize$002,
  input  logic [   0:0] decode_child_serialize$003,
  input  logic [   0:0] decode_child_serialize$004,
  input  logic [   0:0] decode_child_serialize$005,
  input  logic [   0:0] decode_child_serialize$006,
  input  logic [   0:0] decode_child_speculative$000,
  input  logic [   0:0] decode_child_speculative$001,
  input  logic [   0:0] decode_child_speculative$002,
  input  logic [   0:0] decode_child_speculative$003,
  input  logic [   0:0] decode_child_speculative$004,
  input  logic [   0:0] decode_child_speculative$005,
  input  logic [   0:0] decode_child_speculative$006,
  input  logic [   0:0] decode_child_success$000,
  input  logic [   0:0] decode_child_success$001,
  input  logic [   0:0] decode_child_success$002,
  input  logic [   0:0] decode_child_success$003,
  input  logic [   0:0] decode_child_success$004,
  input  logic [   0:0] decode_child_success$005,
  input  logic [   0:0] decode_child_success$006,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // rest_decoder temporaries
  logic   [   0:0] rest_decoder$decode_child_serialize$000;
  logic   [   0:0] rest_decoder$decode_child_serialize$001;
  logic   [   0:0] rest_decoder$decode_child_serialize$002;
  logic   [   0:0] rest_decoder$decode_child_serialize$003;
  logic   [   0:0] rest_decoder$decode_child_serialize$004;
  logic   [   0:0] rest_decoder$decode_child_serialize$005;
  logic   [  14:0] rest_decoder$decode_child_result$000;
  logic   [  14:0] rest_decoder$decode_child_result$001;
  logic   [  14:0] rest_decoder$decode_child_result$002;
  logic   [  14:0] rest_decoder$decode_child_result$003;
  logic   [  14:0] rest_decoder$decode_child_result$004;
  logic   [  14:0] rest_decoder$decode_child_result$005;
  logic   [   0:0] rest_decoder$decode_child_imm_val$000;
  logic   [   0:0] rest_decoder$decode_child_imm_val$001;
  logic   [   0:0] rest_decoder$decode_child_imm_val$002;
  logic   [   0:0] rest_decoder$decode_child_imm_val$003;
  logic   [   0:0] rest_decoder$decode_child_imm_val$004;
  logic   [   0:0] rest_decoder$decode_child_imm_val$005;
  logic   [   0:0] rest_decoder$clk;
  logic   [   2:0] rest_decoder$decode_child_op_class$000;
  logic   [   2:0] rest_decoder$decode_child_op_class$001;
  logic   [   2:0] rest_decoder$decode_child_op_class$002;
  logic   [   2:0] rest_decoder$decode_child_op_class$003;
  logic   [   2:0] rest_decoder$decode_child_op_class$004;
  logic   [   2:0] rest_decoder$decode_child_op_class$005;
  logic   [  31:0] rest_decoder$decode_inst;
  logic   [   0:0] rest_decoder$decode_child_rd_val$000;
  logic   [   0:0] rest_decoder$decode_child_rd_val$001;
  logic   [   0:0] rest_decoder$decode_child_rd_val$002;
  logic   [   0:0] rest_decoder$decode_child_rd_val$003;
  logic   [   0:0] rest_decoder$decode_child_rd_val$004;
  logic   [   0:0] rest_decoder$decode_child_rd_val$005;
  logic   [   0:0] rest_decoder$decode_child_speculative$000;
  logic   [   0:0] rest_decoder$decode_child_speculative$001;
  logic   [   0:0] rest_decoder$decode_child_speculative$002;
  logic   [   0:0] rest_decoder$decode_child_speculative$003;
  logic   [   0:0] rest_decoder$decode_child_speculative$004;
  logic   [   0:0] rest_decoder$decode_child_speculative$005;
  logic   [   0:0] rest_decoder$decode_child_success$000;
  logic   [   0:0] rest_decoder$decode_child_success$001;
  logic   [   0:0] rest_decoder$decode_child_success$002;
  logic   [   0:0] rest_decoder$decode_child_success$003;
  logic   [   0:0] rest_decoder$decode_child_success$004;
  logic   [   0:0] rest_decoder$decode_child_success$005;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$000;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$001;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$002;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$003;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$004;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$005;
  logic   [   0:0] rest_decoder$reset;
  logic   [   2:0] rest_decoder$decode_child_imm_type$000;
  logic   [   2:0] rest_decoder$decode_child_imm_type$001;
  logic   [   2:0] rest_decoder$decode_child_imm_type$002;
  logic   [   2:0] rest_decoder$decode_child_imm_type$003;
  logic   [   2:0] rest_decoder$decode_child_imm_type$004;
  logic   [   2:0] rest_decoder$decode_child_imm_type$005;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$000;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$001;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$002;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$003;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$004;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$005;
  logic   [   2:0] rest_decoder$decode_imm_type;
  logic   [  31:0] rest_decoder$decode_child_inst$000;
  logic   [  31:0] rest_decoder$decode_child_inst$001;
  logic   [  31:0] rest_decoder$decode_child_inst$002;
  logic   [  31:0] rest_decoder$decode_child_inst$003;
  logic   [  31:0] rest_decoder$decode_child_inst$004;
  logic   [  31:0] rest_decoder$decode_child_inst$005;
  logic   [   0:0] rest_decoder$decode_serialize;
  logic   [  14:0] rest_decoder$decode_result;
  logic   [   0:0] rest_decoder$decode_imm_val;
  logic   [   0:0] rest_decoder$decode_rd_val;
  logic   [   0:0] rest_decoder$decode_rs2_val;
  logic   [   2:0] rest_decoder$decode_op_class;
  logic   [   0:0] rest_decoder$decode_success;
  logic   [   0:0] rest_decoder$decode_speculative;
  logic   [   0:0] rest_decoder$decode_rs1_val;

  CompositeDecoder_0x2c27817f255b6f7d rest_decoder
  (
    .decode_child_serialize$000   ( rest_decoder$decode_child_serialize$000 ),
    .decode_child_serialize$001   ( rest_decoder$decode_child_serialize$001 ),
    .decode_child_serialize$002   ( rest_decoder$decode_child_serialize$002 ),
    .decode_child_serialize$003   ( rest_decoder$decode_child_serialize$003 ),
    .decode_child_serialize$004   ( rest_decoder$decode_child_serialize$004 ),
    .decode_child_serialize$005   ( rest_decoder$decode_child_serialize$005 ),
    .decode_child_result$000      ( rest_decoder$decode_child_result$000 ),
    .decode_child_result$001      ( rest_decoder$decode_child_result$001 ),
    .decode_child_result$002      ( rest_decoder$decode_child_result$002 ),
    .decode_child_result$003      ( rest_decoder$decode_child_result$003 ),
    .decode_child_result$004      ( rest_decoder$decode_child_result$004 ),
    .decode_child_result$005      ( rest_decoder$decode_child_result$005 ),
    .decode_child_imm_val$000     ( rest_decoder$decode_child_imm_val$000 ),
    .decode_child_imm_val$001     ( rest_decoder$decode_child_imm_val$001 ),
    .decode_child_imm_val$002     ( rest_decoder$decode_child_imm_val$002 ),
    .decode_child_imm_val$003     ( rest_decoder$decode_child_imm_val$003 ),
    .decode_child_imm_val$004     ( rest_decoder$decode_child_imm_val$004 ),
    .decode_child_imm_val$005     ( rest_decoder$decode_child_imm_val$005 ),
    .clk                          ( rest_decoder$clk ),
    .decode_child_op_class$000    ( rest_decoder$decode_child_op_class$000 ),
    .decode_child_op_class$001    ( rest_decoder$decode_child_op_class$001 ),
    .decode_child_op_class$002    ( rest_decoder$decode_child_op_class$002 ),
    .decode_child_op_class$003    ( rest_decoder$decode_child_op_class$003 ),
    .decode_child_op_class$004    ( rest_decoder$decode_child_op_class$004 ),
    .decode_child_op_class$005    ( rest_decoder$decode_child_op_class$005 ),
    .decode_inst                  ( rest_decoder$decode_inst ),
    .decode_child_rd_val$000      ( rest_decoder$decode_child_rd_val$000 ),
    .decode_child_rd_val$001      ( rest_decoder$decode_child_rd_val$001 ),
    .decode_child_rd_val$002      ( rest_decoder$decode_child_rd_val$002 ),
    .decode_child_rd_val$003      ( rest_decoder$decode_child_rd_val$003 ),
    .decode_child_rd_val$004      ( rest_decoder$decode_child_rd_val$004 ),
    .decode_child_rd_val$005      ( rest_decoder$decode_child_rd_val$005 ),
    .decode_child_speculative$000 ( rest_decoder$decode_child_speculative$000 ),
    .decode_child_speculative$001 ( rest_decoder$decode_child_speculative$001 ),
    .decode_child_speculative$002 ( rest_decoder$decode_child_speculative$002 ),
    .decode_child_speculative$003 ( rest_decoder$decode_child_speculative$003 ),
    .decode_child_speculative$004 ( rest_decoder$decode_child_speculative$004 ),
    .decode_child_speculative$005 ( rest_decoder$decode_child_speculative$005 ),
    .decode_child_success$000     ( rest_decoder$decode_child_success$000 ),
    .decode_child_success$001     ( rest_decoder$decode_child_success$001 ),
    .decode_child_success$002     ( rest_decoder$decode_child_success$002 ),
    .decode_child_success$003     ( rest_decoder$decode_child_success$003 ),
    .decode_child_success$004     ( rest_decoder$decode_child_success$004 ),
    .decode_child_success$005     ( rest_decoder$decode_child_success$005 ),
    .decode_child_rs2_val$000     ( rest_decoder$decode_child_rs2_val$000 ),
    .decode_child_rs2_val$001     ( rest_decoder$decode_child_rs2_val$001 ),
    .decode_child_rs2_val$002     ( rest_decoder$decode_child_rs2_val$002 ),
    .decode_child_rs2_val$003     ( rest_decoder$decode_child_rs2_val$003 ),
    .decode_child_rs2_val$004     ( rest_decoder$decode_child_rs2_val$004 ),
    .decode_child_rs2_val$005     ( rest_decoder$decode_child_rs2_val$005 ),
    .reset                        ( rest_decoder$reset ),
    .decode_child_imm_type$000    ( rest_decoder$decode_child_imm_type$000 ),
    .decode_child_imm_type$001    ( rest_decoder$decode_child_imm_type$001 ),
    .decode_child_imm_type$002    ( rest_decoder$decode_child_imm_type$002 ),
    .decode_child_imm_type$003    ( rest_decoder$decode_child_imm_type$003 ),
    .decode_child_imm_type$004    ( rest_decoder$decode_child_imm_type$004 ),
    .decode_child_imm_type$005    ( rest_decoder$decode_child_imm_type$005 ),
    .decode_child_rs1_val$000     ( rest_decoder$decode_child_rs1_val$000 ),
    .decode_child_rs1_val$001     ( rest_decoder$decode_child_rs1_val$001 ),
    .decode_child_rs1_val$002     ( rest_decoder$decode_child_rs1_val$002 ),
    .decode_child_rs1_val$003     ( rest_decoder$decode_child_rs1_val$003 ),
    .decode_child_rs1_val$004     ( rest_decoder$decode_child_rs1_val$004 ),
    .decode_child_rs1_val$005     ( rest_decoder$decode_child_rs1_val$005 ),
    .decode_imm_type              ( rest_decoder$decode_imm_type ),
    .decode_child_inst$000        ( rest_decoder$decode_child_inst$000 ),
    .decode_child_inst$001        ( rest_decoder$decode_child_inst$001 ),
    .decode_child_inst$002        ( rest_decoder$decode_child_inst$002 ),
    .decode_child_inst$003        ( rest_decoder$decode_child_inst$003 ),
    .decode_child_inst$004        ( rest_decoder$decode_child_inst$004 ),
    .decode_child_inst$005        ( rest_decoder$decode_child_inst$005 ),
    .decode_serialize             ( rest_decoder$decode_serialize ),
    .decode_result                ( rest_decoder$decode_result ),
    .decode_imm_val               ( rest_decoder$decode_imm_val ),
    .decode_rd_val                ( rest_decoder$decode_rd_val ),
    .decode_rs2_val               ( rest_decoder$decode_rs2_val ),
    .decode_op_class              ( rest_decoder$decode_op_class ),
    .decode_success               ( rest_decoder$decode_success ),
    .decode_speculative           ( rest_decoder$decode_speculative ),
    .decode_rs1_val               ( rest_decoder$decode_rs1_val )
  );

  // binary_decoder temporaries
  logic   [   0:0] binary_decoder$decode_b_rs1_val;
  logic   [   0:0] binary_decoder$decode_a_rs1_val;
  logic   [   0:0] binary_decoder$decode_b_rs2_val;
  logic   [   0:0] binary_decoder$decode_a_serialize;
  logic   [  14:0] binary_decoder$decode_a_result;
  logic   [   0:0] binary_decoder$clk;
  logic   [   2:0] binary_decoder$decode_a_imm_type;
  logic   [  31:0] binary_decoder$decode_inst;
  logic   [   0:0] binary_decoder$decode_b_rd_val;
  logic   [   0:0] binary_decoder$decode_a_speculative;
  logic   [   0:0] binary_decoder$decode_a_imm_val;
  logic   [   0:0] binary_decoder$decode_b_success;
  logic   [   2:0] binary_decoder$decode_a_op_class;
  logic   [   0:0] binary_decoder$reset;
  logic   [   2:0] binary_decoder$decode_b_op_class;
  logic   [   2:0] binary_decoder$decode_b_imm_type;
  logic   [   0:0] binary_decoder$decode_a_rd_val;
  logic   [   0:0] binary_decoder$decode_a_success;
  logic   [   0:0] binary_decoder$decode_b_serialize;
  logic   [   0:0] binary_decoder$decode_b_speculative;
  logic   [  14:0] binary_decoder$decode_b_result;
  logic   [   0:0] binary_decoder$decode_a_rs2_val;
  logic   [   0:0] binary_decoder$decode_b_imm_val;
  logic   [   2:0] binary_decoder$decode_imm_type;
  logic   [  31:0] binary_decoder$decode_a_inst;
  logic   [   0:0] binary_decoder$decode_serialize;
  logic   [  14:0] binary_decoder$decode_result;
  logic   [   0:0] binary_decoder$decode_imm_val;
  logic   [   0:0] binary_decoder$decode_rd_val;
  logic   [   0:0] binary_decoder$decode_rs2_val;
  logic   [   2:0] binary_decoder$decode_op_class;
  logic   [   0:0] binary_decoder$decode_success;
  logic   [   0:0] binary_decoder$decode_speculative;
  logic   [  31:0] binary_decoder$decode_b_inst;
  logic   [   0:0] binary_decoder$decode_rs1_val;

  BinaryCompositeDecoder_0x6047cbf454b06e40 binary_decoder
  (
    .decode_b_rs1_val     ( binary_decoder$decode_b_rs1_val ),
    .decode_a_rs1_val     ( binary_decoder$decode_a_rs1_val ),
    .decode_b_rs2_val     ( binary_decoder$decode_b_rs2_val ),
    .decode_a_serialize   ( binary_decoder$decode_a_serialize ),
    .decode_a_result      ( binary_decoder$decode_a_result ),
    .clk                  ( binary_decoder$clk ),
    .decode_a_imm_type    ( binary_decoder$decode_a_imm_type ),
    .decode_inst          ( binary_decoder$decode_inst ),
    .decode_b_rd_val      ( binary_decoder$decode_b_rd_val ),
    .decode_a_speculative ( binary_decoder$decode_a_speculative ),
    .decode_a_imm_val     ( binary_decoder$decode_a_imm_val ),
    .decode_b_success     ( binary_decoder$decode_b_success ),
    .decode_a_op_class    ( binary_decoder$decode_a_op_class ),
    .reset                ( binary_decoder$reset ),
    .decode_b_op_class    ( binary_decoder$decode_b_op_class ),
    .decode_b_imm_type    ( binary_decoder$decode_b_imm_type ),
    .decode_a_rd_val      ( binary_decoder$decode_a_rd_val ),
    .decode_a_success     ( binary_decoder$decode_a_success ),
    .decode_b_serialize   ( binary_decoder$decode_b_serialize ),
    .decode_b_speculative ( binary_decoder$decode_b_speculative ),
    .decode_b_result      ( binary_decoder$decode_b_result ),
    .decode_a_rs2_val     ( binary_decoder$decode_a_rs2_val ),
    .decode_b_imm_val     ( binary_decoder$decode_b_imm_val ),
    .decode_imm_type      ( binary_decoder$decode_imm_type ),
    .decode_a_inst        ( binary_decoder$decode_a_inst ),
    .decode_serialize     ( binary_decoder$decode_serialize ),
    .decode_result        ( binary_decoder$decode_result ),
    .decode_imm_val       ( binary_decoder$decode_imm_val ),
    .decode_rd_val        ( binary_decoder$decode_rd_val ),
    .decode_rs2_val       ( binary_decoder$decode_rs2_val ),
    .decode_op_class      ( binary_decoder$decode_op_class ),
    .decode_success       ( binary_decoder$decode_success ),
    .decode_speculative   ( binary_decoder$decode_speculative ),
    .decode_b_inst        ( binary_decoder$decode_b_inst ),
    .decode_rs1_val       ( binary_decoder$decode_rs1_val )
  );

  // signal connections
  assign binary_decoder$clk                        = clk;
  assign binary_decoder$decode_a_imm_type          = decode_child_imm_type$000;
  assign binary_decoder$decode_a_imm_val           = decode_child_imm_val$000;
  assign binary_decoder$decode_a_op_class          = decode_child_op_class$000;
  assign binary_decoder$decode_a_rd_val            = decode_child_rd_val$000;
  assign binary_decoder$decode_a_result            = decode_child_result$000;
  assign binary_decoder$decode_a_rs1_val           = decode_child_rs1_val$000;
  assign binary_decoder$decode_a_rs2_val           = decode_child_rs2_val$000;
  assign binary_decoder$decode_a_serialize         = decode_child_serialize$000;
  assign binary_decoder$decode_a_speculative       = decode_child_speculative$000;
  assign binary_decoder$decode_a_success           = decode_child_success$000;
  assign binary_decoder$decode_b_imm_type          = rest_decoder$decode_imm_type;
  assign binary_decoder$decode_b_imm_val           = rest_decoder$decode_imm_val;
  assign binary_decoder$decode_b_op_class          = rest_decoder$decode_op_class;
  assign binary_decoder$decode_b_rd_val            = rest_decoder$decode_rd_val;
  assign binary_decoder$decode_b_result            = rest_decoder$decode_result;
  assign binary_decoder$decode_b_rs1_val           = rest_decoder$decode_rs1_val;
  assign binary_decoder$decode_b_rs2_val           = rest_decoder$decode_rs2_val;
  assign binary_decoder$decode_b_serialize         = rest_decoder$decode_serialize;
  assign binary_decoder$decode_b_speculative       = rest_decoder$decode_speculative;
  assign binary_decoder$decode_b_success           = rest_decoder$decode_success;
  assign binary_decoder$decode_inst                = decode_inst;
  assign binary_decoder$reset                      = reset;
  assign decode_child_inst$000                     = binary_decoder$decode_a_inst;
  assign decode_child_inst$001                     = rest_decoder$decode_child_inst$000;
  assign decode_child_inst$002                     = rest_decoder$decode_child_inst$001;
  assign decode_child_inst$003                     = rest_decoder$decode_child_inst$002;
  assign decode_child_inst$004                     = rest_decoder$decode_child_inst$003;
  assign decode_child_inst$005                     = rest_decoder$decode_child_inst$004;
  assign decode_child_inst$006                     = rest_decoder$decode_child_inst$005;
  assign decode_imm_type                           = binary_decoder$decode_imm_type;
  assign decode_imm_val                            = binary_decoder$decode_imm_val;
  assign decode_op_class                           = binary_decoder$decode_op_class;
  assign decode_rd_val                             = binary_decoder$decode_rd_val;
  assign decode_result                             = binary_decoder$decode_result;
  assign decode_rs1_val                            = binary_decoder$decode_rs1_val;
  assign decode_rs2_val                            = binary_decoder$decode_rs2_val;
  assign decode_serialize                          = binary_decoder$decode_serialize;
  assign decode_speculative                        = binary_decoder$decode_speculative;
  assign decode_success                            = binary_decoder$decode_success;
  assign rest_decoder$clk                          = clk;
  assign rest_decoder$decode_child_imm_type$000    = decode_child_imm_type$001;
  assign rest_decoder$decode_child_imm_type$001    = decode_child_imm_type$002;
  assign rest_decoder$decode_child_imm_type$002    = decode_child_imm_type$003;
  assign rest_decoder$decode_child_imm_type$003    = decode_child_imm_type$004;
  assign rest_decoder$decode_child_imm_type$004    = decode_child_imm_type$005;
  assign rest_decoder$decode_child_imm_type$005    = decode_child_imm_type$006;
  assign rest_decoder$decode_child_imm_val$000     = decode_child_imm_val$001;
  assign rest_decoder$decode_child_imm_val$001     = decode_child_imm_val$002;
  assign rest_decoder$decode_child_imm_val$002     = decode_child_imm_val$003;
  assign rest_decoder$decode_child_imm_val$003     = decode_child_imm_val$004;
  assign rest_decoder$decode_child_imm_val$004     = decode_child_imm_val$005;
  assign rest_decoder$decode_child_imm_val$005     = decode_child_imm_val$006;
  assign rest_decoder$decode_child_op_class$000    = decode_child_op_class$001;
  assign rest_decoder$decode_child_op_class$001    = decode_child_op_class$002;
  assign rest_decoder$decode_child_op_class$002    = decode_child_op_class$003;
  assign rest_decoder$decode_child_op_class$003    = decode_child_op_class$004;
  assign rest_decoder$decode_child_op_class$004    = decode_child_op_class$005;
  assign rest_decoder$decode_child_op_class$005    = decode_child_op_class$006;
  assign rest_decoder$decode_child_rd_val$000      = decode_child_rd_val$001;
  assign rest_decoder$decode_child_rd_val$001      = decode_child_rd_val$002;
  assign rest_decoder$decode_child_rd_val$002      = decode_child_rd_val$003;
  assign rest_decoder$decode_child_rd_val$003      = decode_child_rd_val$004;
  assign rest_decoder$decode_child_rd_val$004      = decode_child_rd_val$005;
  assign rest_decoder$decode_child_rd_val$005      = decode_child_rd_val$006;
  assign rest_decoder$decode_child_result$000      = decode_child_result$001;
  assign rest_decoder$decode_child_result$001      = decode_child_result$002;
  assign rest_decoder$decode_child_result$002      = decode_child_result$003;
  assign rest_decoder$decode_child_result$003      = decode_child_result$004;
  assign rest_decoder$decode_child_result$004      = decode_child_result$005;
  assign rest_decoder$decode_child_result$005      = decode_child_result$006;
  assign rest_decoder$decode_child_rs1_val$000     = decode_child_rs1_val$001;
  assign rest_decoder$decode_child_rs1_val$001     = decode_child_rs1_val$002;
  assign rest_decoder$decode_child_rs1_val$002     = decode_child_rs1_val$003;
  assign rest_decoder$decode_child_rs1_val$003     = decode_child_rs1_val$004;
  assign rest_decoder$decode_child_rs1_val$004     = decode_child_rs1_val$005;
  assign rest_decoder$decode_child_rs1_val$005     = decode_child_rs1_val$006;
  assign rest_decoder$decode_child_rs2_val$000     = decode_child_rs2_val$001;
  assign rest_decoder$decode_child_rs2_val$001     = decode_child_rs2_val$002;
  assign rest_decoder$decode_child_rs2_val$002     = decode_child_rs2_val$003;
  assign rest_decoder$decode_child_rs2_val$003     = decode_child_rs2_val$004;
  assign rest_decoder$decode_child_rs2_val$004     = decode_child_rs2_val$005;
  assign rest_decoder$decode_child_rs2_val$005     = decode_child_rs2_val$006;
  assign rest_decoder$decode_child_serialize$000   = decode_child_serialize$001;
  assign rest_decoder$decode_child_serialize$001   = decode_child_serialize$002;
  assign rest_decoder$decode_child_serialize$002   = decode_child_serialize$003;
  assign rest_decoder$decode_child_serialize$003   = decode_child_serialize$004;
  assign rest_decoder$decode_child_serialize$004   = decode_child_serialize$005;
  assign rest_decoder$decode_child_serialize$005   = decode_child_serialize$006;
  assign rest_decoder$decode_child_speculative$000 = decode_child_speculative$001;
  assign rest_decoder$decode_child_speculative$001 = decode_child_speculative$002;
  assign rest_decoder$decode_child_speculative$002 = decode_child_speculative$003;
  assign rest_decoder$decode_child_speculative$003 = decode_child_speculative$004;
  assign rest_decoder$decode_child_speculative$004 = decode_child_speculative$005;
  assign rest_decoder$decode_child_speculative$005 = decode_child_speculative$006;
  assign rest_decoder$decode_child_success$000     = decode_child_success$001;
  assign rest_decoder$decode_child_success$001     = decode_child_success$002;
  assign rest_decoder$decode_child_success$002     = decode_child_success$003;
  assign rest_decoder$decode_child_success$003     = decode_child_success$004;
  assign rest_decoder$decode_child_success$004     = decode_child_success$005;
  assign rest_decoder$decode_child_success$005     = decode_child_success$006;
  assign rest_decoder$decode_inst                  = binary_decoder$decode_b_inst;
  assign rest_decoder$reset                        = reset;



endmodule // CompositeDecoder_0x2c27817f254c2cc0

//-----------------------------------------------------------------------------
// CompositeDecoder_0x2c27817f255b6f7d
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"nchildren": 6}
// PyMTL: verilator_xinit = zeros
module CompositeDecoder_0x2c27817f255b6f7d
(
  input  logic [   0:0] clk,
  input  logic [   2:0] decode_child_imm_type$000,
  input  logic [   2:0] decode_child_imm_type$001,
  input  logic [   2:0] decode_child_imm_type$002,
  input  logic [   2:0] decode_child_imm_type$003,
  input  logic [   2:0] decode_child_imm_type$004,
  input  logic [   2:0] decode_child_imm_type$005,
  input  logic [   0:0] decode_child_imm_val$000,
  input  logic [   0:0] decode_child_imm_val$001,
  input  logic [   0:0] decode_child_imm_val$002,
  input  logic [   0:0] decode_child_imm_val$003,
  input  logic [   0:0] decode_child_imm_val$004,
  input  logic [   0:0] decode_child_imm_val$005,
  output logic [  31:0] decode_child_inst$000,
  output logic [  31:0] decode_child_inst$001,
  output logic [  31:0] decode_child_inst$002,
  output logic [  31:0] decode_child_inst$003,
  output logic [  31:0] decode_child_inst$004,
  output logic [  31:0] decode_child_inst$005,
  input  logic [   2:0] decode_child_op_class$000,
  input  logic [   2:0] decode_child_op_class$001,
  input  logic [   2:0] decode_child_op_class$002,
  input  logic [   2:0] decode_child_op_class$003,
  input  logic [   2:0] decode_child_op_class$004,
  input  logic [   2:0] decode_child_op_class$005,
  input  logic [   0:0] decode_child_rd_val$000,
  input  logic [   0:0] decode_child_rd_val$001,
  input  logic [   0:0] decode_child_rd_val$002,
  input  logic [   0:0] decode_child_rd_val$003,
  input  logic [   0:0] decode_child_rd_val$004,
  input  logic [   0:0] decode_child_rd_val$005,
  input  logic [  14:0] decode_child_result$000,
  input  logic [  14:0] decode_child_result$001,
  input  logic [  14:0] decode_child_result$002,
  input  logic [  14:0] decode_child_result$003,
  input  logic [  14:0] decode_child_result$004,
  input  logic [  14:0] decode_child_result$005,
  input  logic [   0:0] decode_child_rs1_val$000,
  input  logic [   0:0] decode_child_rs1_val$001,
  input  logic [   0:0] decode_child_rs1_val$002,
  input  logic [   0:0] decode_child_rs1_val$003,
  input  logic [   0:0] decode_child_rs1_val$004,
  input  logic [   0:0] decode_child_rs1_val$005,
  input  logic [   0:0] decode_child_rs2_val$000,
  input  logic [   0:0] decode_child_rs2_val$001,
  input  logic [   0:0] decode_child_rs2_val$002,
  input  logic [   0:0] decode_child_rs2_val$003,
  input  logic [   0:0] decode_child_rs2_val$004,
  input  logic [   0:0] decode_child_rs2_val$005,
  input  logic [   0:0] decode_child_serialize$000,
  input  logic [   0:0] decode_child_serialize$001,
  input  logic [   0:0] decode_child_serialize$002,
  input  logic [   0:0] decode_child_serialize$003,
  input  logic [   0:0] decode_child_serialize$004,
  input  logic [   0:0] decode_child_serialize$005,
  input  logic [   0:0] decode_child_speculative$000,
  input  logic [   0:0] decode_child_speculative$001,
  input  logic [   0:0] decode_child_speculative$002,
  input  logic [   0:0] decode_child_speculative$003,
  input  logic [   0:0] decode_child_speculative$004,
  input  logic [   0:0] decode_child_speculative$005,
  input  logic [   0:0] decode_child_success$000,
  input  logic [   0:0] decode_child_success$001,
  input  logic [   0:0] decode_child_success$002,
  input  logic [   0:0] decode_child_success$003,
  input  logic [   0:0] decode_child_success$004,
  input  logic [   0:0] decode_child_success$005,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // rest_decoder temporaries
  logic   [   0:0] rest_decoder$decode_child_serialize$000;
  logic   [   0:0] rest_decoder$decode_child_serialize$001;
  logic   [   0:0] rest_decoder$decode_child_serialize$002;
  logic   [   0:0] rest_decoder$decode_child_serialize$003;
  logic   [   0:0] rest_decoder$decode_child_serialize$004;
  logic   [  14:0] rest_decoder$decode_child_result$000;
  logic   [  14:0] rest_decoder$decode_child_result$001;
  logic   [  14:0] rest_decoder$decode_child_result$002;
  logic   [  14:0] rest_decoder$decode_child_result$003;
  logic   [  14:0] rest_decoder$decode_child_result$004;
  logic   [   0:0] rest_decoder$decode_child_imm_val$000;
  logic   [   0:0] rest_decoder$decode_child_imm_val$001;
  logic   [   0:0] rest_decoder$decode_child_imm_val$002;
  logic   [   0:0] rest_decoder$decode_child_imm_val$003;
  logic   [   0:0] rest_decoder$decode_child_imm_val$004;
  logic   [   0:0] rest_decoder$clk;
  logic   [   2:0] rest_decoder$decode_child_op_class$000;
  logic   [   2:0] rest_decoder$decode_child_op_class$001;
  logic   [   2:0] rest_decoder$decode_child_op_class$002;
  logic   [   2:0] rest_decoder$decode_child_op_class$003;
  logic   [   2:0] rest_decoder$decode_child_op_class$004;
  logic   [  31:0] rest_decoder$decode_inst;
  logic   [   0:0] rest_decoder$decode_child_rd_val$000;
  logic   [   0:0] rest_decoder$decode_child_rd_val$001;
  logic   [   0:0] rest_decoder$decode_child_rd_val$002;
  logic   [   0:0] rest_decoder$decode_child_rd_val$003;
  logic   [   0:0] rest_decoder$decode_child_rd_val$004;
  logic   [   0:0] rest_decoder$decode_child_speculative$000;
  logic   [   0:0] rest_decoder$decode_child_speculative$001;
  logic   [   0:0] rest_decoder$decode_child_speculative$002;
  logic   [   0:0] rest_decoder$decode_child_speculative$003;
  logic   [   0:0] rest_decoder$decode_child_speculative$004;
  logic   [   0:0] rest_decoder$decode_child_success$000;
  logic   [   0:0] rest_decoder$decode_child_success$001;
  logic   [   0:0] rest_decoder$decode_child_success$002;
  logic   [   0:0] rest_decoder$decode_child_success$003;
  logic   [   0:0] rest_decoder$decode_child_success$004;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$000;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$001;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$002;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$003;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$004;
  logic   [   0:0] rest_decoder$reset;
  logic   [   2:0] rest_decoder$decode_child_imm_type$000;
  logic   [   2:0] rest_decoder$decode_child_imm_type$001;
  logic   [   2:0] rest_decoder$decode_child_imm_type$002;
  logic   [   2:0] rest_decoder$decode_child_imm_type$003;
  logic   [   2:0] rest_decoder$decode_child_imm_type$004;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$000;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$001;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$002;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$003;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$004;
  logic   [   2:0] rest_decoder$decode_imm_type;
  logic   [  31:0] rest_decoder$decode_child_inst$000;
  logic   [  31:0] rest_decoder$decode_child_inst$001;
  logic   [  31:0] rest_decoder$decode_child_inst$002;
  logic   [  31:0] rest_decoder$decode_child_inst$003;
  logic   [  31:0] rest_decoder$decode_child_inst$004;
  logic   [   0:0] rest_decoder$decode_serialize;
  logic   [  14:0] rest_decoder$decode_result;
  logic   [   0:0] rest_decoder$decode_imm_val;
  logic   [   0:0] rest_decoder$decode_rd_val;
  logic   [   0:0] rest_decoder$decode_rs2_val;
  logic   [   2:0] rest_decoder$decode_op_class;
  logic   [   0:0] rest_decoder$decode_success;
  logic   [   0:0] rest_decoder$decode_speculative;
  logic   [   0:0] rest_decoder$decode_rs1_val;

  CompositeDecoder_0x2c27817f252da836 rest_decoder
  (
    .decode_child_serialize$000   ( rest_decoder$decode_child_serialize$000 ),
    .decode_child_serialize$001   ( rest_decoder$decode_child_serialize$001 ),
    .decode_child_serialize$002   ( rest_decoder$decode_child_serialize$002 ),
    .decode_child_serialize$003   ( rest_decoder$decode_child_serialize$003 ),
    .decode_child_serialize$004   ( rest_decoder$decode_child_serialize$004 ),
    .decode_child_result$000      ( rest_decoder$decode_child_result$000 ),
    .decode_child_result$001      ( rest_decoder$decode_child_result$001 ),
    .decode_child_result$002      ( rest_decoder$decode_child_result$002 ),
    .decode_child_result$003      ( rest_decoder$decode_child_result$003 ),
    .decode_child_result$004      ( rest_decoder$decode_child_result$004 ),
    .decode_child_imm_val$000     ( rest_decoder$decode_child_imm_val$000 ),
    .decode_child_imm_val$001     ( rest_decoder$decode_child_imm_val$001 ),
    .decode_child_imm_val$002     ( rest_decoder$decode_child_imm_val$002 ),
    .decode_child_imm_val$003     ( rest_decoder$decode_child_imm_val$003 ),
    .decode_child_imm_val$004     ( rest_decoder$decode_child_imm_val$004 ),
    .clk                          ( rest_decoder$clk ),
    .decode_child_op_class$000    ( rest_decoder$decode_child_op_class$000 ),
    .decode_child_op_class$001    ( rest_decoder$decode_child_op_class$001 ),
    .decode_child_op_class$002    ( rest_decoder$decode_child_op_class$002 ),
    .decode_child_op_class$003    ( rest_decoder$decode_child_op_class$003 ),
    .decode_child_op_class$004    ( rest_decoder$decode_child_op_class$004 ),
    .decode_inst                  ( rest_decoder$decode_inst ),
    .decode_child_rd_val$000      ( rest_decoder$decode_child_rd_val$000 ),
    .decode_child_rd_val$001      ( rest_decoder$decode_child_rd_val$001 ),
    .decode_child_rd_val$002      ( rest_decoder$decode_child_rd_val$002 ),
    .decode_child_rd_val$003      ( rest_decoder$decode_child_rd_val$003 ),
    .decode_child_rd_val$004      ( rest_decoder$decode_child_rd_val$004 ),
    .decode_child_speculative$000 ( rest_decoder$decode_child_speculative$000 ),
    .decode_child_speculative$001 ( rest_decoder$decode_child_speculative$001 ),
    .decode_child_speculative$002 ( rest_decoder$decode_child_speculative$002 ),
    .decode_child_speculative$003 ( rest_decoder$decode_child_speculative$003 ),
    .decode_child_speculative$004 ( rest_decoder$decode_child_speculative$004 ),
    .decode_child_success$000     ( rest_decoder$decode_child_success$000 ),
    .decode_child_success$001     ( rest_decoder$decode_child_success$001 ),
    .decode_child_success$002     ( rest_decoder$decode_child_success$002 ),
    .decode_child_success$003     ( rest_decoder$decode_child_success$003 ),
    .decode_child_success$004     ( rest_decoder$decode_child_success$004 ),
    .decode_child_rs2_val$000     ( rest_decoder$decode_child_rs2_val$000 ),
    .decode_child_rs2_val$001     ( rest_decoder$decode_child_rs2_val$001 ),
    .decode_child_rs2_val$002     ( rest_decoder$decode_child_rs2_val$002 ),
    .decode_child_rs2_val$003     ( rest_decoder$decode_child_rs2_val$003 ),
    .decode_child_rs2_val$004     ( rest_decoder$decode_child_rs2_val$004 ),
    .reset                        ( rest_decoder$reset ),
    .decode_child_imm_type$000    ( rest_decoder$decode_child_imm_type$000 ),
    .decode_child_imm_type$001    ( rest_decoder$decode_child_imm_type$001 ),
    .decode_child_imm_type$002    ( rest_decoder$decode_child_imm_type$002 ),
    .decode_child_imm_type$003    ( rest_decoder$decode_child_imm_type$003 ),
    .decode_child_imm_type$004    ( rest_decoder$decode_child_imm_type$004 ),
    .decode_child_rs1_val$000     ( rest_decoder$decode_child_rs1_val$000 ),
    .decode_child_rs1_val$001     ( rest_decoder$decode_child_rs1_val$001 ),
    .decode_child_rs1_val$002     ( rest_decoder$decode_child_rs1_val$002 ),
    .decode_child_rs1_val$003     ( rest_decoder$decode_child_rs1_val$003 ),
    .decode_child_rs1_val$004     ( rest_decoder$decode_child_rs1_val$004 ),
    .decode_imm_type              ( rest_decoder$decode_imm_type ),
    .decode_child_inst$000        ( rest_decoder$decode_child_inst$000 ),
    .decode_child_inst$001        ( rest_decoder$decode_child_inst$001 ),
    .decode_child_inst$002        ( rest_decoder$decode_child_inst$002 ),
    .decode_child_inst$003        ( rest_decoder$decode_child_inst$003 ),
    .decode_child_inst$004        ( rest_decoder$decode_child_inst$004 ),
    .decode_serialize             ( rest_decoder$decode_serialize ),
    .decode_result                ( rest_decoder$decode_result ),
    .decode_imm_val               ( rest_decoder$decode_imm_val ),
    .decode_rd_val                ( rest_decoder$decode_rd_val ),
    .decode_rs2_val               ( rest_decoder$decode_rs2_val ),
    .decode_op_class              ( rest_decoder$decode_op_class ),
    .decode_success               ( rest_decoder$decode_success ),
    .decode_speculative           ( rest_decoder$decode_speculative ),
    .decode_rs1_val               ( rest_decoder$decode_rs1_val )
  );

  // binary_decoder temporaries
  logic   [   0:0] binary_decoder$decode_b_rs1_val;
  logic   [   0:0] binary_decoder$decode_a_rs1_val;
  logic   [   0:0] binary_decoder$decode_b_rs2_val;
  logic   [   0:0] binary_decoder$decode_a_serialize;
  logic   [  14:0] binary_decoder$decode_a_result;
  logic   [   0:0] binary_decoder$clk;
  logic   [   2:0] binary_decoder$decode_a_imm_type;
  logic   [  31:0] binary_decoder$decode_inst;
  logic   [   0:0] binary_decoder$decode_b_rd_val;
  logic   [   0:0] binary_decoder$decode_a_speculative;
  logic   [   0:0] binary_decoder$decode_a_imm_val;
  logic   [   0:0] binary_decoder$decode_b_success;
  logic   [   2:0] binary_decoder$decode_a_op_class;
  logic   [   0:0] binary_decoder$reset;
  logic   [   2:0] binary_decoder$decode_b_op_class;
  logic   [   2:0] binary_decoder$decode_b_imm_type;
  logic   [   0:0] binary_decoder$decode_a_rd_val;
  logic   [   0:0] binary_decoder$decode_a_success;
  logic   [   0:0] binary_decoder$decode_b_serialize;
  logic   [   0:0] binary_decoder$decode_b_speculative;
  logic   [  14:0] binary_decoder$decode_b_result;
  logic   [   0:0] binary_decoder$decode_a_rs2_val;
  logic   [   0:0] binary_decoder$decode_b_imm_val;
  logic   [   2:0] binary_decoder$decode_imm_type;
  logic   [  31:0] binary_decoder$decode_a_inst;
  logic   [   0:0] binary_decoder$decode_serialize;
  logic   [  14:0] binary_decoder$decode_result;
  logic   [   0:0] binary_decoder$decode_imm_val;
  logic   [   0:0] binary_decoder$decode_rd_val;
  logic   [   0:0] binary_decoder$decode_rs2_val;
  logic   [   2:0] binary_decoder$decode_op_class;
  logic   [   0:0] binary_decoder$decode_success;
  logic   [   0:0] binary_decoder$decode_speculative;
  logic   [  31:0] binary_decoder$decode_b_inst;
  logic   [   0:0] binary_decoder$decode_rs1_val;

  BinaryCompositeDecoder_0x6047cbf454b06e40 binary_decoder
  (
    .decode_b_rs1_val     ( binary_decoder$decode_b_rs1_val ),
    .decode_a_rs1_val     ( binary_decoder$decode_a_rs1_val ),
    .decode_b_rs2_val     ( binary_decoder$decode_b_rs2_val ),
    .decode_a_serialize   ( binary_decoder$decode_a_serialize ),
    .decode_a_result      ( binary_decoder$decode_a_result ),
    .clk                  ( binary_decoder$clk ),
    .decode_a_imm_type    ( binary_decoder$decode_a_imm_type ),
    .decode_inst          ( binary_decoder$decode_inst ),
    .decode_b_rd_val      ( binary_decoder$decode_b_rd_val ),
    .decode_a_speculative ( binary_decoder$decode_a_speculative ),
    .decode_a_imm_val     ( binary_decoder$decode_a_imm_val ),
    .decode_b_success     ( binary_decoder$decode_b_success ),
    .decode_a_op_class    ( binary_decoder$decode_a_op_class ),
    .reset                ( binary_decoder$reset ),
    .decode_b_op_class    ( binary_decoder$decode_b_op_class ),
    .decode_b_imm_type    ( binary_decoder$decode_b_imm_type ),
    .decode_a_rd_val      ( binary_decoder$decode_a_rd_val ),
    .decode_a_success     ( binary_decoder$decode_a_success ),
    .decode_b_serialize   ( binary_decoder$decode_b_serialize ),
    .decode_b_speculative ( binary_decoder$decode_b_speculative ),
    .decode_b_result      ( binary_decoder$decode_b_result ),
    .decode_a_rs2_val     ( binary_decoder$decode_a_rs2_val ),
    .decode_b_imm_val     ( binary_decoder$decode_b_imm_val ),
    .decode_imm_type      ( binary_decoder$decode_imm_type ),
    .decode_a_inst        ( binary_decoder$decode_a_inst ),
    .decode_serialize     ( binary_decoder$decode_serialize ),
    .decode_result        ( binary_decoder$decode_result ),
    .decode_imm_val       ( binary_decoder$decode_imm_val ),
    .decode_rd_val        ( binary_decoder$decode_rd_val ),
    .decode_rs2_val       ( binary_decoder$decode_rs2_val ),
    .decode_op_class      ( binary_decoder$decode_op_class ),
    .decode_success       ( binary_decoder$decode_success ),
    .decode_speculative   ( binary_decoder$decode_speculative ),
    .decode_b_inst        ( binary_decoder$decode_b_inst ),
    .decode_rs1_val       ( binary_decoder$decode_rs1_val )
  );

  // signal connections
  assign binary_decoder$clk                        = clk;
  assign binary_decoder$decode_a_imm_type          = decode_child_imm_type$000;
  assign binary_decoder$decode_a_imm_val           = decode_child_imm_val$000;
  assign binary_decoder$decode_a_op_class          = decode_child_op_class$000;
  assign binary_decoder$decode_a_rd_val            = decode_child_rd_val$000;
  assign binary_decoder$decode_a_result            = decode_child_result$000;
  assign binary_decoder$decode_a_rs1_val           = decode_child_rs1_val$000;
  assign binary_decoder$decode_a_rs2_val           = decode_child_rs2_val$000;
  assign binary_decoder$decode_a_serialize         = decode_child_serialize$000;
  assign binary_decoder$decode_a_speculative       = decode_child_speculative$000;
  assign binary_decoder$decode_a_success           = decode_child_success$000;
  assign binary_decoder$decode_b_imm_type          = rest_decoder$decode_imm_type;
  assign binary_decoder$decode_b_imm_val           = rest_decoder$decode_imm_val;
  assign binary_decoder$decode_b_op_class          = rest_decoder$decode_op_class;
  assign binary_decoder$decode_b_rd_val            = rest_decoder$decode_rd_val;
  assign binary_decoder$decode_b_result            = rest_decoder$decode_result;
  assign binary_decoder$decode_b_rs1_val           = rest_decoder$decode_rs1_val;
  assign binary_decoder$decode_b_rs2_val           = rest_decoder$decode_rs2_val;
  assign binary_decoder$decode_b_serialize         = rest_decoder$decode_serialize;
  assign binary_decoder$decode_b_speculative       = rest_decoder$decode_speculative;
  assign binary_decoder$decode_b_success           = rest_decoder$decode_success;
  assign binary_decoder$decode_inst                = decode_inst;
  assign binary_decoder$reset                      = reset;
  assign decode_child_inst$000                     = binary_decoder$decode_a_inst;
  assign decode_child_inst$001                     = rest_decoder$decode_child_inst$000;
  assign decode_child_inst$002                     = rest_decoder$decode_child_inst$001;
  assign decode_child_inst$003                     = rest_decoder$decode_child_inst$002;
  assign decode_child_inst$004                     = rest_decoder$decode_child_inst$003;
  assign decode_child_inst$005                     = rest_decoder$decode_child_inst$004;
  assign decode_imm_type                           = binary_decoder$decode_imm_type;
  assign decode_imm_val                            = binary_decoder$decode_imm_val;
  assign decode_op_class                           = binary_decoder$decode_op_class;
  assign decode_rd_val                             = binary_decoder$decode_rd_val;
  assign decode_result                             = binary_decoder$decode_result;
  assign decode_rs1_val                            = binary_decoder$decode_rs1_val;
  assign decode_rs2_val                            = binary_decoder$decode_rs2_val;
  assign decode_serialize                          = binary_decoder$decode_serialize;
  assign decode_speculative                        = binary_decoder$decode_speculative;
  assign decode_success                            = binary_decoder$decode_success;
  assign rest_decoder$clk                          = clk;
  assign rest_decoder$decode_child_imm_type$000    = decode_child_imm_type$001;
  assign rest_decoder$decode_child_imm_type$001    = decode_child_imm_type$002;
  assign rest_decoder$decode_child_imm_type$002    = decode_child_imm_type$003;
  assign rest_decoder$decode_child_imm_type$003    = decode_child_imm_type$004;
  assign rest_decoder$decode_child_imm_type$004    = decode_child_imm_type$005;
  assign rest_decoder$decode_child_imm_val$000     = decode_child_imm_val$001;
  assign rest_decoder$decode_child_imm_val$001     = decode_child_imm_val$002;
  assign rest_decoder$decode_child_imm_val$002     = decode_child_imm_val$003;
  assign rest_decoder$decode_child_imm_val$003     = decode_child_imm_val$004;
  assign rest_decoder$decode_child_imm_val$004     = decode_child_imm_val$005;
  assign rest_decoder$decode_child_op_class$000    = decode_child_op_class$001;
  assign rest_decoder$decode_child_op_class$001    = decode_child_op_class$002;
  assign rest_decoder$decode_child_op_class$002    = decode_child_op_class$003;
  assign rest_decoder$decode_child_op_class$003    = decode_child_op_class$004;
  assign rest_decoder$decode_child_op_class$004    = decode_child_op_class$005;
  assign rest_decoder$decode_child_rd_val$000      = decode_child_rd_val$001;
  assign rest_decoder$decode_child_rd_val$001      = decode_child_rd_val$002;
  assign rest_decoder$decode_child_rd_val$002      = decode_child_rd_val$003;
  assign rest_decoder$decode_child_rd_val$003      = decode_child_rd_val$004;
  assign rest_decoder$decode_child_rd_val$004      = decode_child_rd_val$005;
  assign rest_decoder$decode_child_result$000      = decode_child_result$001;
  assign rest_decoder$decode_child_result$001      = decode_child_result$002;
  assign rest_decoder$decode_child_result$002      = decode_child_result$003;
  assign rest_decoder$decode_child_result$003      = decode_child_result$004;
  assign rest_decoder$decode_child_result$004      = decode_child_result$005;
  assign rest_decoder$decode_child_rs1_val$000     = decode_child_rs1_val$001;
  assign rest_decoder$decode_child_rs1_val$001     = decode_child_rs1_val$002;
  assign rest_decoder$decode_child_rs1_val$002     = decode_child_rs1_val$003;
  assign rest_decoder$decode_child_rs1_val$003     = decode_child_rs1_val$004;
  assign rest_decoder$decode_child_rs1_val$004     = decode_child_rs1_val$005;
  assign rest_decoder$decode_child_rs2_val$000     = decode_child_rs2_val$001;
  assign rest_decoder$decode_child_rs2_val$001     = decode_child_rs2_val$002;
  assign rest_decoder$decode_child_rs2_val$002     = decode_child_rs2_val$003;
  assign rest_decoder$decode_child_rs2_val$003     = decode_child_rs2_val$004;
  assign rest_decoder$decode_child_rs2_val$004     = decode_child_rs2_val$005;
  assign rest_decoder$decode_child_serialize$000   = decode_child_serialize$001;
  assign rest_decoder$decode_child_serialize$001   = decode_child_serialize$002;
  assign rest_decoder$decode_child_serialize$002   = decode_child_serialize$003;
  assign rest_decoder$decode_child_serialize$003   = decode_child_serialize$004;
  assign rest_decoder$decode_child_serialize$004   = decode_child_serialize$005;
  assign rest_decoder$decode_child_speculative$000 = decode_child_speculative$001;
  assign rest_decoder$decode_child_speculative$001 = decode_child_speculative$002;
  assign rest_decoder$decode_child_speculative$002 = decode_child_speculative$003;
  assign rest_decoder$decode_child_speculative$003 = decode_child_speculative$004;
  assign rest_decoder$decode_child_speculative$004 = decode_child_speculative$005;
  assign rest_decoder$decode_child_success$000     = decode_child_success$001;
  assign rest_decoder$decode_child_success$001     = decode_child_success$002;
  assign rest_decoder$decode_child_success$002     = decode_child_success$003;
  assign rest_decoder$decode_child_success$003     = decode_child_success$004;
  assign rest_decoder$decode_child_success$004     = decode_child_success$005;
  assign rest_decoder$decode_inst                  = binary_decoder$decode_b_inst;
  assign rest_decoder$reset                        = reset;



endmodule // CompositeDecoder_0x2c27817f255b6f7d

//-----------------------------------------------------------------------------
// CompositeDecoder_0x2c27817f252da836
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"nchildren": 5}
// PyMTL: verilator_xinit = zeros
module CompositeDecoder_0x2c27817f252da836
(
  input  logic [   0:0] clk,
  input  logic [   2:0] decode_child_imm_type$000,
  input  logic [   2:0] decode_child_imm_type$001,
  input  logic [   2:0] decode_child_imm_type$002,
  input  logic [   2:0] decode_child_imm_type$003,
  input  logic [   2:0] decode_child_imm_type$004,
  input  logic [   0:0] decode_child_imm_val$000,
  input  logic [   0:0] decode_child_imm_val$001,
  input  logic [   0:0] decode_child_imm_val$002,
  input  logic [   0:0] decode_child_imm_val$003,
  input  logic [   0:0] decode_child_imm_val$004,
  output logic [  31:0] decode_child_inst$000,
  output logic [  31:0] decode_child_inst$001,
  output logic [  31:0] decode_child_inst$002,
  output logic [  31:0] decode_child_inst$003,
  output logic [  31:0] decode_child_inst$004,
  input  logic [   2:0] decode_child_op_class$000,
  input  logic [   2:0] decode_child_op_class$001,
  input  logic [   2:0] decode_child_op_class$002,
  input  logic [   2:0] decode_child_op_class$003,
  input  logic [   2:0] decode_child_op_class$004,
  input  logic [   0:0] decode_child_rd_val$000,
  input  logic [   0:0] decode_child_rd_val$001,
  input  logic [   0:0] decode_child_rd_val$002,
  input  logic [   0:0] decode_child_rd_val$003,
  input  logic [   0:0] decode_child_rd_val$004,
  input  logic [  14:0] decode_child_result$000,
  input  logic [  14:0] decode_child_result$001,
  input  logic [  14:0] decode_child_result$002,
  input  logic [  14:0] decode_child_result$003,
  input  logic [  14:0] decode_child_result$004,
  input  logic [   0:0] decode_child_rs1_val$000,
  input  logic [   0:0] decode_child_rs1_val$001,
  input  logic [   0:0] decode_child_rs1_val$002,
  input  logic [   0:0] decode_child_rs1_val$003,
  input  logic [   0:0] decode_child_rs1_val$004,
  input  logic [   0:0] decode_child_rs2_val$000,
  input  logic [   0:0] decode_child_rs2_val$001,
  input  logic [   0:0] decode_child_rs2_val$002,
  input  logic [   0:0] decode_child_rs2_val$003,
  input  logic [   0:0] decode_child_rs2_val$004,
  input  logic [   0:0] decode_child_serialize$000,
  input  logic [   0:0] decode_child_serialize$001,
  input  logic [   0:0] decode_child_serialize$002,
  input  logic [   0:0] decode_child_serialize$003,
  input  logic [   0:0] decode_child_serialize$004,
  input  logic [   0:0] decode_child_speculative$000,
  input  logic [   0:0] decode_child_speculative$001,
  input  logic [   0:0] decode_child_speculative$002,
  input  logic [   0:0] decode_child_speculative$003,
  input  logic [   0:0] decode_child_speculative$004,
  input  logic [   0:0] decode_child_success$000,
  input  logic [   0:0] decode_child_success$001,
  input  logic [   0:0] decode_child_success$002,
  input  logic [   0:0] decode_child_success$003,
  input  logic [   0:0] decode_child_success$004,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // rest_decoder temporaries
  logic   [   0:0] rest_decoder$decode_child_serialize$000;
  logic   [   0:0] rest_decoder$decode_child_serialize$001;
  logic   [   0:0] rest_decoder$decode_child_serialize$002;
  logic   [   0:0] rest_decoder$decode_child_serialize$003;
  logic   [  14:0] rest_decoder$decode_child_result$000;
  logic   [  14:0] rest_decoder$decode_child_result$001;
  logic   [  14:0] rest_decoder$decode_child_result$002;
  logic   [  14:0] rest_decoder$decode_child_result$003;
  logic   [   0:0] rest_decoder$decode_child_imm_val$000;
  logic   [   0:0] rest_decoder$decode_child_imm_val$001;
  logic   [   0:0] rest_decoder$decode_child_imm_val$002;
  logic   [   0:0] rest_decoder$decode_child_imm_val$003;
  logic   [   0:0] rest_decoder$clk;
  logic   [   2:0] rest_decoder$decode_child_op_class$000;
  logic   [   2:0] rest_decoder$decode_child_op_class$001;
  logic   [   2:0] rest_decoder$decode_child_op_class$002;
  logic   [   2:0] rest_decoder$decode_child_op_class$003;
  logic   [  31:0] rest_decoder$decode_inst;
  logic   [   0:0] rest_decoder$decode_child_rd_val$000;
  logic   [   0:0] rest_decoder$decode_child_rd_val$001;
  logic   [   0:0] rest_decoder$decode_child_rd_val$002;
  logic   [   0:0] rest_decoder$decode_child_rd_val$003;
  logic   [   0:0] rest_decoder$decode_child_speculative$000;
  logic   [   0:0] rest_decoder$decode_child_speculative$001;
  logic   [   0:0] rest_decoder$decode_child_speculative$002;
  logic   [   0:0] rest_decoder$decode_child_speculative$003;
  logic   [   0:0] rest_decoder$decode_child_success$000;
  logic   [   0:0] rest_decoder$decode_child_success$001;
  logic   [   0:0] rest_decoder$decode_child_success$002;
  logic   [   0:0] rest_decoder$decode_child_success$003;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$000;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$001;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$002;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$003;
  logic   [   0:0] rest_decoder$reset;
  logic   [   2:0] rest_decoder$decode_child_imm_type$000;
  logic   [   2:0] rest_decoder$decode_child_imm_type$001;
  logic   [   2:0] rest_decoder$decode_child_imm_type$002;
  logic   [   2:0] rest_decoder$decode_child_imm_type$003;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$000;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$001;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$002;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$003;
  logic   [   2:0] rest_decoder$decode_imm_type;
  logic   [  31:0] rest_decoder$decode_child_inst$000;
  logic   [  31:0] rest_decoder$decode_child_inst$001;
  logic   [  31:0] rest_decoder$decode_child_inst$002;
  logic   [  31:0] rest_decoder$decode_child_inst$003;
  logic   [   0:0] rest_decoder$decode_serialize;
  logic   [  14:0] rest_decoder$decode_result;
  logic   [   0:0] rest_decoder$decode_imm_val;
  logic   [   0:0] rest_decoder$decode_rd_val;
  logic   [   0:0] rest_decoder$decode_rs2_val;
  logic   [   2:0] rest_decoder$decode_op_class;
  logic   [   0:0] rest_decoder$decode_success;
  logic   [   0:0] rest_decoder$decode_speculative;
  logic   [   0:0] rest_decoder$decode_rs1_val;

  CompositeDecoder_0x2c27817f253ceafb rest_decoder
  (
    .decode_child_serialize$000   ( rest_decoder$decode_child_serialize$000 ),
    .decode_child_serialize$001   ( rest_decoder$decode_child_serialize$001 ),
    .decode_child_serialize$002   ( rest_decoder$decode_child_serialize$002 ),
    .decode_child_serialize$003   ( rest_decoder$decode_child_serialize$003 ),
    .decode_child_result$000      ( rest_decoder$decode_child_result$000 ),
    .decode_child_result$001      ( rest_decoder$decode_child_result$001 ),
    .decode_child_result$002      ( rest_decoder$decode_child_result$002 ),
    .decode_child_result$003      ( rest_decoder$decode_child_result$003 ),
    .decode_child_imm_val$000     ( rest_decoder$decode_child_imm_val$000 ),
    .decode_child_imm_val$001     ( rest_decoder$decode_child_imm_val$001 ),
    .decode_child_imm_val$002     ( rest_decoder$decode_child_imm_val$002 ),
    .decode_child_imm_val$003     ( rest_decoder$decode_child_imm_val$003 ),
    .clk                          ( rest_decoder$clk ),
    .decode_child_op_class$000    ( rest_decoder$decode_child_op_class$000 ),
    .decode_child_op_class$001    ( rest_decoder$decode_child_op_class$001 ),
    .decode_child_op_class$002    ( rest_decoder$decode_child_op_class$002 ),
    .decode_child_op_class$003    ( rest_decoder$decode_child_op_class$003 ),
    .decode_inst                  ( rest_decoder$decode_inst ),
    .decode_child_rd_val$000      ( rest_decoder$decode_child_rd_val$000 ),
    .decode_child_rd_val$001      ( rest_decoder$decode_child_rd_val$001 ),
    .decode_child_rd_val$002      ( rest_decoder$decode_child_rd_val$002 ),
    .decode_child_rd_val$003      ( rest_decoder$decode_child_rd_val$003 ),
    .decode_child_speculative$000 ( rest_decoder$decode_child_speculative$000 ),
    .decode_child_speculative$001 ( rest_decoder$decode_child_speculative$001 ),
    .decode_child_speculative$002 ( rest_decoder$decode_child_speculative$002 ),
    .decode_child_speculative$003 ( rest_decoder$decode_child_speculative$003 ),
    .decode_child_success$000     ( rest_decoder$decode_child_success$000 ),
    .decode_child_success$001     ( rest_decoder$decode_child_success$001 ),
    .decode_child_success$002     ( rest_decoder$decode_child_success$002 ),
    .decode_child_success$003     ( rest_decoder$decode_child_success$003 ),
    .decode_child_rs2_val$000     ( rest_decoder$decode_child_rs2_val$000 ),
    .decode_child_rs2_val$001     ( rest_decoder$decode_child_rs2_val$001 ),
    .decode_child_rs2_val$002     ( rest_decoder$decode_child_rs2_val$002 ),
    .decode_child_rs2_val$003     ( rest_decoder$decode_child_rs2_val$003 ),
    .reset                        ( rest_decoder$reset ),
    .decode_child_imm_type$000    ( rest_decoder$decode_child_imm_type$000 ),
    .decode_child_imm_type$001    ( rest_decoder$decode_child_imm_type$001 ),
    .decode_child_imm_type$002    ( rest_decoder$decode_child_imm_type$002 ),
    .decode_child_imm_type$003    ( rest_decoder$decode_child_imm_type$003 ),
    .decode_child_rs1_val$000     ( rest_decoder$decode_child_rs1_val$000 ),
    .decode_child_rs1_val$001     ( rest_decoder$decode_child_rs1_val$001 ),
    .decode_child_rs1_val$002     ( rest_decoder$decode_child_rs1_val$002 ),
    .decode_child_rs1_val$003     ( rest_decoder$decode_child_rs1_val$003 ),
    .decode_imm_type              ( rest_decoder$decode_imm_type ),
    .decode_child_inst$000        ( rest_decoder$decode_child_inst$000 ),
    .decode_child_inst$001        ( rest_decoder$decode_child_inst$001 ),
    .decode_child_inst$002        ( rest_decoder$decode_child_inst$002 ),
    .decode_child_inst$003        ( rest_decoder$decode_child_inst$003 ),
    .decode_serialize             ( rest_decoder$decode_serialize ),
    .decode_result                ( rest_decoder$decode_result ),
    .decode_imm_val               ( rest_decoder$decode_imm_val ),
    .decode_rd_val                ( rest_decoder$decode_rd_val ),
    .decode_rs2_val               ( rest_decoder$decode_rs2_val ),
    .decode_op_class              ( rest_decoder$decode_op_class ),
    .decode_success               ( rest_decoder$decode_success ),
    .decode_speculative           ( rest_decoder$decode_speculative ),
    .decode_rs1_val               ( rest_decoder$decode_rs1_val )
  );

  // binary_decoder temporaries
  logic   [   0:0] binary_decoder$decode_b_rs1_val;
  logic   [   0:0] binary_decoder$decode_a_rs1_val;
  logic   [   0:0] binary_decoder$decode_b_rs2_val;
  logic   [   0:0] binary_decoder$decode_a_serialize;
  logic   [  14:0] binary_decoder$decode_a_result;
  logic   [   0:0] binary_decoder$clk;
  logic   [   2:0] binary_decoder$decode_a_imm_type;
  logic   [  31:0] binary_decoder$decode_inst;
  logic   [   0:0] binary_decoder$decode_b_rd_val;
  logic   [   0:0] binary_decoder$decode_a_speculative;
  logic   [   0:0] binary_decoder$decode_a_imm_val;
  logic   [   0:0] binary_decoder$decode_b_success;
  logic   [   2:0] binary_decoder$decode_a_op_class;
  logic   [   0:0] binary_decoder$reset;
  logic   [   2:0] binary_decoder$decode_b_op_class;
  logic   [   2:0] binary_decoder$decode_b_imm_type;
  logic   [   0:0] binary_decoder$decode_a_rd_val;
  logic   [   0:0] binary_decoder$decode_a_success;
  logic   [   0:0] binary_decoder$decode_b_serialize;
  logic   [   0:0] binary_decoder$decode_b_speculative;
  logic   [  14:0] binary_decoder$decode_b_result;
  logic   [   0:0] binary_decoder$decode_a_rs2_val;
  logic   [   0:0] binary_decoder$decode_b_imm_val;
  logic   [   2:0] binary_decoder$decode_imm_type;
  logic   [  31:0] binary_decoder$decode_a_inst;
  logic   [   0:0] binary_decoder$decode_serialize;
  logic   [  14:0] binary_decoder$decode_result;
  logic   [   0:0] binary_decoder$decode_imm_val;
  logic   [   0:0] binary_decoder$decode_rd_val;
  logic   [   0:0] binary_decoder$decode_rs2_val;
  logic   [   2:0] binary_decoder$decode_op_class;
  logic   [   0:0] binary_decoder$decode_success;
  logic   [   0:0] binary_decoder$decode_speculative;
  logic   [  31:0] binary_decoder$decode_b_inst;
  logic   [   0:0] binary_decoder$decode_rs1_val;

  BinaryCompositeDecoder_0x6047cbf454b06e40 binary_decoder
  (
    .decode_b_rs1_val     ( binary_decoder$decode_b_rs1_val ),
    .decode_a_rs1_val     ( binary_decoder$decode_a_rs1_val ),
    .decode_b_rs2_val     ( binary_decoder$decode_b_rs2_val ),
    .decode_a_serialize   ( binary_decoder$decode_a_serialize ),
    .decode_a_result      ( binary_decoder$decode_a_result ),
    .clk                  ( binary_decoder$clk ),
    .decode_a_imm_type    ( binary_decoder$decode_a_imm_type ),
    .decode_inst          ( binary_decoder$decode_inst ),
    .decode_b_rd_val      ( binary_decoder$decode_b_rd_val ),
    .decode_a_speculative ( binary_decoder$decode_a_speculative ),
    .decode_a_imm_val     ( binary_decoder$decode_a_imm_val ),
    .decode_b_success     ( binary_decoder$decode_b_success ),
    .decode_a_op_class    ( binary_decoder$decode_a_op_class ),
    .reset                ( binary_decoder$reset ),
    .decode_b_op_class    ( binary_decoder$decode_b_op_class ),
    .decode_b_imm_type    ( binary_decoder$decode_b_imm_type ),
    .decode_a_rd_val      ( binary_decoder$decode_a_rd_val ),
    .decode_a_success     ( binary_decoder$decode_a_success ),
    .decode_b_serialize   ( binary_decoder$decode_b_serialize ),
    .decode_b_speculative ( binary_decoder$decode_b_speculative ),
    .decode_b_result      ( binary_decoder$decode_b_result ),
    .decode_a_rs2_val     ( binary_decoder$decode_a_rs2_val ),
    .decode_b_imm_val     ( binary_decoder$decode_b_imm_val ),
    .decode_imm_type      ( binary_decoder$decode_imm_type ),
    .decode_a_inst        ( binary_decoder$decode_a_inst ),
    .decode_serialize     ( binary_decoder$decode_serialize ),
    .decode_result        ( binary_decoder$decode_result ),
    .decode_imm_val       ( binary_decoder$decode_imm_val ),
    .decode_rd_val        ( binary_decoder$decode_rd_val ),
    .decode_rs2_val       ( binary_decoder$decode_rs2_val ),
    .decode_op_class      ( binary_decoder$decode_op_class ),
    .decode_success       ( binary_decoder$decode_success ),
    .decode_speculative   ( binary_decoder$decode_speculative ),
    .decode_b_inst        ( binary_decoder$decode_b_inst ),
    .decode_rs1_val       ( binary_decoder$decode_rs1_val )
  );

  // signal connections
  assign binary_decoder$clk                        = clk;
  assign binary_decoder$decode_a_imm_type          = decode_child_imm_type$000;
  assign binary_decoder$decode_a_imm_val           = decode_child_imm_val$000;
  assign binary_decoder$decode_a_op_class          = decode_child_op_class$000;
  assign binary_decoder$decode_a_rd_val            = decode_child_rd_val$000;
  assign binary_decoder$decode_a_result            = decode_child_result$000;
  assign binary_decoder$decode_a_rs1_val           = decode_child_rs1_val$000;
  assign binary_decoder$decode_a_rs2_val           = decode_child_rs2_val$000;
  assign binary_decoder$decode_a_serialize         = decode_child_serialize$000;
  assign binary_decoder$decode_a_speculative       = decode_child_speculative$000;
  assign binary_decoder$decode_a_success           = decode_child_success$000;
  assign binary_decoder$decode_b_imm_type          = rest_decoder$decode_imm_type;
  assign binary_decoder$decode_b_imm_val           = rest_decoder$decode_imm_val;
  assign binary_decoder$decode_b_op_class          = rest_decoder$decode_op_class;
  assign binary_decoder$decode_b_rd_val            = rest_decoder$decode_rd_val;
  assign binary_decoder$decode_b_result            = rest_decoder$decode_result;
  assign binary_decoder$decode_b_rs1_val           = rest_decoder$decode_rs1_val;
  assign binary_decoder$decode_b_rs2_val           = rest_decoder$decode_rs2_val;
  assign binary_decoder$decode_b_serialize         = rest_decoder$decode_serialize;
  assign binary_decoder$decode_b_speculative       = rest_decoder$decode_speculative;
  assign binary_decoder$decode_b_success           = rest_decoder$decode_success;
  assign binary_decoder$decode_inst                = decode_inst;
  assign binary_decoder$reset                      = reset;
  assign decode_child_inst$000                     = binary_decoder$decode_a_inst;
  assign decode_child_inst$001                     = rest_decoder$decode_child_inst$000;
  assign decode_child_inst$002                     = rest_decoder$decode_child_inst$001;
  assign decode_child_inst$003                     = rest_decoder$decode_child_inst$002;
  assign decode_child_inst$004                     = rest_decoder$decode_child_inst$003;
  assign decode_imm_type                           = binary_decoder$decode_imm_type;
  assign decode_imm_val                            = binary_decoder$decode_imm_val;
  assign decode_op_class                           = binary_decoder$decode_op_class;
  assign decode_rd_val                             = binary_decoder$decode_rd_val;
  assign decode_result                             = binary_decoder$decode_result;
  assign decode_rs1_val                            = binary_decoder$decode_rs1_val;
  assign decode_rs2_val                            = binary_decoder$decode_rs2_val;
  assign decode_serialize                          = binary_decoder$decode_serialize;
  assign decode_speculative                        = binary_decoder$decode_speculative;
  assign decode_success                            = binary_decoder$decode_success;
  assign rest_decoder$clk                          = clk;
  assign rest_decoder$decode_child_imm_type$000    = decode_child_imm_type$001;
  assign rest_decoder$decode_child_imm_type$001    = decode_child_imm_type$002;
  assign rest_decoder$decode_child_imm_type$002    = decode_child_imm_type$003;
  assign rest_decoder$decode_child_imm_type$003    = decode_child_imm_type$004;
  assign rest_decoder$decode_child_imm_val$000     = decode_child_imm_val$001;
  assign rest_decoder$decode_child_imm_val$001     = decode_child_imm_val$002;
  assign rest_decoder$decode_child_imm_val$002     = decode_child_imm_val$003;
  assign rest_decoder$decode_child_imm_val$003     = decode_child_imm_val$004;
  assign rest_decoder$decode_child_op_class$000    = decode_child_op_class$001;
  assign rest_decoder$decode_child_op_class$001    = decode_child_op_class$002;
  assign rest_decoder$decode_child_op_class$002    = decode_child_op_class$003;
  assign rest_decoder$decode_child_op_class$003    = decode_child_op_class$004;
  assign rest_decoder$decode_child_rd_val$000      = decode_child_rd_val$001;
  assign rest_decoder$decode_child_rd_val$001      = decode_child_rd_val$002;
  assign rest_decoder$decode_child_rd_val$002      = decode_child_rd_val$003;
  assign rest_decoder$decode_child_rd_val$003      = decode_child_rd_val$004;
  assign rest_decoder$decode_child_result$000      = decode_child_result$001;
  assign rest_decoder$decode_child_result$001      = decode_child_result$002;
  assign rest_decoder$decode_child_result$002      = decode_child_result$003;
  assign rest_decoder$decode_child_result$003      = decode_child_result$004;
  assign rest_decoder$decode_child_rs1_val$000     = decode_child_rs1_val$001;
  assign rest_decoder$decode_child_rs1_val$001     = decode_child_rs1_val$002;
  assign rest_decoder$decode_child_rs1_val$002     = decode_child_rs1_val$003;
  assign rest_decoder$decode_child_rs1_val$003     = decode_child_rs1_val$004;
  assign rest_decoder$decode_child_rs2_val$000     = decode_child_rs2_val$001;
  assign rest_decoder$decode_child_rs2_val$001     = decode_child_rs2_val$002;
  assign rest_decoder$decode_child_rs2_val$002     = decode_child_rs2_val$003;
  assign rest_decoder$decode_child_rs2_val$003     = decode_child_rs2_val$004;
  assign rest_decoder$decode_child_serialize$000   = decode_child_serialize$001;
  assign rest_decoder$decode_child_serialize$001   = decode_child_serialize$002;
  assign rest_decoder$decode_child_serialize$002   = decode_child_serialize$003;
  assign rest_decoder$decode_child_serialize$003   = decode_child_serialize$004;
  assign rest_decoder$decode_child_speculative$000 = decode_child_speculative$001;
  assign rest_decoder$decode_child_speculative$001 = decode_child_speculative$002;
  assign rest_decoder$decode_child_speculative$002 = decode_child_speculative$003;
  assign rest_decoder$decode_child_speculative$003 = decode_child_speculative$004;
  assign rest_decoder$decode_child_success$000     = decode_child_success$001;
  assign rest_decoder$decode_child_success$001     = decode_child_success$002;
  assign rest_decoder$decode_child_success$002     = decode_child_success$003;
  assign rest_decoder$decode_child_success$003     = decode_child_success$004;
  assign rest_decoder$decode_inst                  = binary_decoder$decode_b_inst;
  assign rest_decoder$reset                        = reset;



endmodule // CompositeDecoder_0x2c27817f252da836

//-----------------------------------------------------------------------------
// CompositeDecoder_0x2c27817f253ceafb
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"nchildren": 4}
// PyMTL: verilator_xinit = zeros
module CompositeDecoder_0x2c27817f253ceafb
(
  input  logic [   0:0] clk,
  input  logic [   2:0] decode_child_imm_type$000,
  input  logic [   2:0] decode_child_imm_type$001,
  input  logic [   2:0] decode_child_imm_type$002,
  input  logic [   2:0] decode_child_imm_type$003,
  input  logic [   0:0] decode_child_imm_val$000,
  input  logic [   0:0] decode_child_imm_val$001,
  input  logic [   0:0] decode_child_imm_val$002,
  input  logic [   0:0] decode_child_imm_val$003,
  output logic [  31:0] decode_child_inst$000,
  output logic [  31:0] decode_child_inst$001,
  output logic [  31:0] decode_child_inst$002,
  output logic [  31:0] decode_child_inst$003,
  input  logic [   2:0] decode_child_op_class$000,
  input  logic [   2:0] decode_child_op_class$001,
  input  logic [   2:0] decode_child_op_class$002,
  input  logic [   2:0] decode_child_op_class$003,
  input  logic [   0:0] decode_child_rd_val$000,
  input  logic [   0:0] decode_child_rd_val$001,
  input  logic [   0:0] decode_child_rd_val$002,
  input  logic [   0:0] decode_child_rd_val$003,
  input  logic [  14:0] decode_child_result$000,
  input  logic [  14:0] decode_child_result$001,
  input  logic [  14:0] decode_child_result$002,
  input  logic [  14:0] decode_child_result$003,
  input  logic [   0:0] decode_child_rs1_val$000,
  input  logic [   0:0] decode_child_rs1_val$001,
  input  logic [   0:0] decode_child_rs1_val$002,
  input  logic [   0:0] decode_child_rs1_val$003,
  input  logic [   0:0] decode_child_rs2_val$000,
  input  logic [   0:0] decode_child_rs2_val$001,
  input  logic [   0:0] decode_child_rs2_val$002,
  input  logic [   0:0] decode_child_rs2_val$003,
  input  logic [   0:0] decode_child_serialize$000,
  input  logic [   0:0] decode_child_serialize$001,
  input  logic [   0:0] decode_child_serialize$002,
  input  logic [   0:0] decode_child_serialize$003,
  input  logic [   0:0] decode_child_speculative$000,
  input  logic [   0:0] decode_child_speculative$001,
  input  logic [   0:0] decode_child_speculative$002,
  input  logic [   0:0] decode_child_speculative$003,
  input  logic [   0:0] decode_child_success$000,
  input  logic [   0:0] decode_child_success$001,
  input  logic [   0:0] decode_child_success$002,
  input  logic [   0:0] decode_child_success$003,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // rest_decoder temporaries
  logic   [   0:0] rest_decoder$decode_child_serialize$000;
  logic   [   0:0] rest_decoder$decode_child_serialize$001;
  logic   [   0:0] rest_decoder$decode_child_serialize$002;
  logic   [  14:0] rest_decoder$decode_child_result$000;
  logic   [  14:0] rest_decoder$decode_child_result$001;
  logic   [  14:0] rest_decoder$decode_child_result$002;
  logic   [   0:0] rest_decoder$decode_child_imm_val$000;
  logic   [   0:0] rest_decoder$decode_child_imm_val$001;
  logic   [   0:0] rest_decoder$decode_child_imm_val$002;
  logic   [   0:0] rest_decoder$clk;
  logic   [   2:0] rest_decoder$decode_child_op_class$000;
  logic   [   2:0] rest_decoder$decode_child_op_class$001;
  logic   [   2:0] rest_decoder$decode_child_op_class$002;
  logic   [  31:0] rest_decoder$decode_inst;
  logic   [   0:0] rest_decoder$decode_child_rd_val$000;
  logic   [   0:0] rest_decoder$decode_child_rd_val$001;
  logic   [   0:0] rest_decoder$decode_child_rd_val$002;
  logic   [   0:0] rest_decoder$decode_child_speculative$000;
  logic   [   0:0] rest_decoder$decode_child_speculative$001;
  logic   [   0:0] rest_decoder$decode_child_speculative$002;
  logic   [   0:0] rest_decoder$decode_child_success$000;
  logic   [   0:0] rest_decoder$decode_child_success$001;
  logic   [   0:0] rest_decoder$decode_child_success$002;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$000;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$001;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$002;
  logic   [   0:0] rest_decoder$reset;
  logic   [   2:0] rest_decoder$decode_child_imm_type$000;
  logic   [   2:0] rest_decoder$decode_child_imm_type$001;
  logic   [   2:0] rest_decoder$decode_child_imm_type$002;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$000;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$001;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$002;
  logic   [   2:0] rest_decoder$decode_imm_type;
  logic   [  31:0] rest_decoder$decode_child_inst$000;
  logic   [  31:0] rest_decoder$decode_child_inst$001;
  logic   [  31:0] rest_decoder$decode_child_inst$002;
  logic   [   0:0] rest_decoder$decode_serialize;
  logic   [  14:0] rest_decoder$decode_result;
  logic   [   0:0] rest_decoder$decode_imm_val;
  logic   [   0:0] rest_decoder$decode_rd_val;
  logic   [   0:0] rest_decoder$decode_rs2_val;
  logic   [   2:0] rest_decoder$decode_op_class;
  logic   [   0:0] rest_decoder$decode_success;
  logic   [   0:0] rest_decoder$decode_speculative;
  logic   [   0:0] rest_decoder$decode_rs1_val;

  CompositeDecoder_0x2c27817f250f23b4 rest_decoder
  (
    .decode_child_serialize$000   ( rest_decoder$decode_child_serialize$000 ),
    .decode_child_serialize$001   ( rest_decoder$decode_child_serialize$001 ),
    .decode_child_serialize$002   ( rest_decoder$decode_child_serialize$002 ),
    .decode_child_result$000      ( rest_decoder$decode_child_result$000 ),
    .decode_child_result$001      ( rest_decoder$decode_child_result$001 ),
    .decode_child_result$002      ( rest_decoder$decode_child_result$002 ),
    .decode_child_imm_val$000     ( rest_decoder$decode_child_imm_val$000 ),
    .decode_child_imm_val$001     ( rest_decoder$decode_child_imm_val$001 ),
    .decode_child_imm_val$002     ( rest_decoder$decode_child_imm_val$002 ),
    .clk                          ( rest_decoder$clk ),
    .decode_child_op_class$000    ( rest_decoder$decode_child_op_class$000 ),
    .decode_child_op_class$001    ( rest_decoder$decode_child_op_class$001 ),
    .decode_child_op_class$002    ( rest_decoder$decode_child_op_class$002 ),
    .decode_inst                  ( rest_decoder$decode_inst ),
    .decode_child_rd_val$000      ( rest_decoder$decode_child_rd_val$000 ),
    .decode_child_rd_val$001      ( rest_decoder$decode_child_rd_val$001 ),
    .decode_child_rd_val$002      ( rest_decoder$decode_child_rd_val$002 ),
    .decode_child_speculative$000 ( rest_decoder$decode_child_speculative$000 ),
    .decode_child_speculative$001 ( rest_decoder$decode_child_speculative$001 ),
    .decode_child_speculative$002 ( rest_decoder$decode_child_speculative$002 ),
    .decode_child_success$000     ( rest_decoder$decode_child_success$000 ),
    .decode_child_success$001     ( rest_decoder$decode_child_success$001 ),
    .decode_child_success$002     ( rest_decoder$decode_child_success$002 ),
    .decode_child_rs2_val$000     ( rest_decoder$decode_child_rs2_val$000 ),
    .decode_child_rs2_val$001     ( rest_decoder$decode_child_rs2_val$001 ),
    .decode_child_rs2_val$002     ( rest_decoder$decode_child_rs2_val$002 ),
    .reset                        ( rest_decoder$reset ),
    .decode_child_imm_type$000    ( rest_decoder$decode_child_imm_type$000 ),
    .decode_child_imm_type$001    ( rest_decoder$decode_child_imm_type$001 ),
    .decode_child_imm_type$002    ( rest_decoder$decode_child_imm_type$002 ),
    .decode_child_rs1_val$000     ( rest_decoder$decode_child_rs1_val$000 ),
    .decode_child_rs1_val$001     ( rest_decoder$decode_child_rs1_val$001 ),
    .decode_child_rs1_val$002     ( rest_decoder$decode_child_rs1_val$002 ),
    .decode_imm_type              ( rest_decoder$decode_imm_type ),
    .decode_child_inst$000        ( rest_decoder$decode_child_inst$000 ),
    .decode_child_inst$001        ( rest_decoder$decode_child_inst$001 ),
    .decode_child_inst$002        ( rest_decoder$decode_child_inst$002 ),
    .decode_serialize             ( rest_decoder$decode_serialize ),
    .decode_result                ( rest_decoder$decode_result ),
    .decode_imm_val               ( rest_decoder$decode_imm_val ),
    .decode_rd_val                ( rest_decoder$decode_rd_val ),
    .decode_rs2_val               ( rest_decoder$decode_rs2_val ),
    .decode_op_class              ( rest_decoder$decode_op_class ),
    .decode_success               ( rest_decoder$decode_success ),
    .decode_speculative           ( rest_decoder$decode_speculative ),
    .decode_rs1_val               ( rest_decoder$decode_rs1_val )
  );

  // binary_decoder temporaries
  logic   [   0:0] binary_decoder$decode_b_rs1_val;
  logic   [   0:0] binary_decoder$decode_a_rs1_val;
  logic   [   0:0] binary_decoder$decode_b_rs2_val;
  logic   [   0:0] binary_decoder$decode_a_serialize;
  logic   [  14:0] binary_decoder$decode_a_result;
  logic   [   0:0] binary_decoder$clk;
  logic   [   2:0] binary_decoder$decode_a_imm_type;
  logic   [  31:0] binary_decoder$decode_inst;
  logic   [   0:0] binary_decoder$decode_b_rd_val;
  logic   [   0:0] binary_decoder$decode_a_speculative;
  logic   [   0:0] binary_decoder$decode_a_imm_val;
  logic   [   0:0] binary_decoder$decode_b_success;
  logic   [   2:0] binary_decoder$decode_a_op_class;
  logic   [   0:0] binary_decoder$reset;
  logic   [   2:0] binary_decoder$decode_b_op_class;
  logic   [   2:0] binary_decoder$decode_b_imm_type;
  logic   [   0:0] binary_decoder$decode_a_rd_val;
  logic   [   0:0] binary_decoder$decode_a_success;
  logic   [   0:0] binary_decoder$decode_b_serialize;
  logic   [   0:0] binary_decoder$decode_b_speculative;
  logic   [  14:0] binary_decoder$decode_b_result;
  logic   [   0:0] binary_decoder$decode_a_rs2_val;
  logic   [   0:0] binary_decoder$decode_b_imm_val;
  logic   [   2:0] binary_decoder$decode_imm_type;
  logic   [  31:0] binary_decoder$decode_a_inst;
  logic   [   0:0] binary_decoder$decode_serialize;
  logic   [  14:0] binary_decoder$decode_result;
  logic   [   0:0] binary_decoder$decode_imm_val;
  logic   [   0:0] binary_decoder$decode_rd_val;
  logic   [   0:0] binary_decoder$decode_rs2_val;
  logic   [   2:0] binary_decoder$decode_op_class;
  logic   [   0:0] binary_decoder$decode_success;
  logic   [   0:0] binary_decoder$decode_speculative;
  logic   [  31:0] binary_decoder$decode_b_inst;
  logic   [   0:0] binary_decoder$decode_rs1_val;

  BinaryCompositeDecoder_0x6047cbf454b06e40 binary_decoder
  (
    .decode_b_rs1_val     ( binary_decoder$decode_b_rs1_val ),
    .decode_a_rs1_val     ( binary_decoder$decode_a_rs1_val ),
    .decode_b_rs2_val     ( binary_decoder$decode_b_rs2_val ),
    .decode_a_serialize   ( binary_decoder$decode_a_serialize ),
    .decode_a_result      ( binary_decoder$decode_a_result ),
    .clk                  ( binary_decoder$clk ),
    .decode_a_imm_type    ( binary_decoder$decode_a_imm_type ),
    .decode_inst          ( binary_decoder$decode_inst ),
    .decode_b_rd_val      ( binary_decoder$decode_b_rd_val ),
    .decode_a_speculative ( binary_decoder$decode_a_speculative ),
    .decode_a_imm_val     ( binary_decoder$decode_a_imm_val ),
    .decode_b_success     ( binary_decoder$decode_b_success ),
    .decode_a_op_class    ( binary_decoder$decode_a_op_class ),
    .reset                ( binary_decoder$reset ),
    .decode_b_op_class    ( binary_decoder$decode_b_op_class ),
    .decode_b_imm_type    ( binary_decoder$decode_b_imm_type ),
    .decode_a_rd_val      ( binary_decoder$decode_a_rd_val ),
    .decode_a_success     ( binary_decoder$decode_a_success ),
    .decode_b_serialize   ( binary_decoder$decode_b_serialize ),
    .decode_b_speculative ( binary_decoder$decode_b_speculative ),
    .decode_b_result      ( binary_decoder$decode_b_result ),
    .decode_a_rs2_val     ( binary_decoder$decode_a_rs2_val ),
    .decode_b_imm_val     ( binary_decoder$decode_b_imm_val ),
    .decode_imm_type      ( binary_decoder$decode_imm_type ),
    .decode_a_inst        ( binary_decoder$decode_a_inst ),
    .decode_serialize     ( binary_decoder$decode_serialize ),
    .decode_result        ( binary_decoder$decode_result ),
    .decode_imm_val       ( binary_decoder$decode_imm_val ),
    .decode_rd_val        ( binary_decoder$decode_rd_val ),
    .decode_rs2_val       ( binary_decoder$decode_rs2_val ),
    .decode_op_class      ( binary_decoder$decode_op_class ),
    .decode_success       ( binary_decoder$decode_success ),
    .decode_speculative   ( binary_decoder$decode_speculative ),
    .decode_b_inst        ( binary_decoder$decode_b_inst ),
    .decode_rs1_val       ( binary_decoder$decode_rs1_val )
  );

  // signal connections
  assign binary_decoder$clk                        = clk;
  assign binary_decoder$decode_a_imm_type          = decode_child_imm_type$000;
  assign binary_decoder$decode_a_imm_val           = decode_child_imm_val$000;
  assign binary_decoder$decode_a_op_class          = decode_child_op_class$000;
  assign binary_decoder$decode_a_rd_val            = decode_child_rd_val$000;
  assign binary_decoder$decode_a_result            = decode_child_result$000;
  assign binary_decoder$decode_a_rs1_val           = decode_child_rs1_val$000;
  assign binary_decoder$decode_a_rs2_val           = decode_child_rs2_val$000;
  assign binary_decoder$decode_a_serialize         = decode_child_serialize$000;
  assign binary_decoder$decode_a_speculative       = decode_child_speculative$000;
  assign binary_decoder$decode_a_success           = decode_child_success$000;
  assign binary_decoder$decode_b_imm_type          = rest_decoder$decode_imm_type;
  assign binary_decoder$decode_b_imm_val           = rest_decoder$decode_imm_val;
  assign binary_decoder$decode_b_op_class          = rest_decoder$decode_op_class;
  assign binary_decoder$decode_b_rd_val            = rest_decoder$decode_rd_val;
  assign binary_decoder$decode_b_result            = rest_decoder$decode_result;
  assign binary_decoder$decode_b_rs1_val           = rest_decoder$decode_rs1_val;
  assign binary_decoder$decode_b_rs2_val           = rest_decoder$decode_rs2_val;
  assign binary_decoder$decode_b_serialize         = rest_decoder$decode_serialize;
  assign binary_decoder$decode_b_speculative       = rest_decoder$decode_speculative;
  assign binary_decoder$decode_b_success           = rest_decoder$decode_success;
  assign binary_decoder$decode_inst                = decode_inst;
  assign binary_decoder$reset                      = reset;
  assign decode_child_inst$000                     = binary_decoder$decode_a_inst;
  assign decode_child_inst$001                     = rest_decoder$decode_child_inst$000;
  assign decode_child_inst$002                     = rest_decoder$decode_child_inst$001;
  assign decode_child_inst$003                     = rest_decoder$decode_child_inst$002;
  assign decode_imm_type                           = binary_decoder$decode_imm_type;
  assign decode_imm_val                            = binary_decoder$decode_imm_val;
  assign decode_op_class                           = binary_decoder$decode_op_class;
  assign decode_rd_val                             = binary_decoder$decode_rd_val;
  assign decode_result                             = binary_decoder$decode_result;
  assign decode_rs1_val                            = binary_decoder$decode_rs1_val;
  assign decode_rs2_val                            = binary_decoder$decode_rs2_val;
  assign decode_serialize                          = binary_decoder$decode_serialize;
  assign decode_speculative                        = binary_decoder$decode_speculative;
  assign decode_success                            = binary_decoder$decode_success;
  assign rest_decoder$clk                          = clk;
  assign rest_decoder$decode_child_imm_type$000    = decode_child_imm_type$001;
  assign rest_decoder$decode_child_imm_type$001    = decode_child_imm_type$002;
  assign rest_decoder$decode_child_imm_type$002    = decode_child_imm_type$003;
  assign rest_decoder$decode_child_imm_val$000     = decode_child_imm_val$001;
  assign rest_decoder$decode_child_imm_val$001     = decode_child_imm_val$002;
  assign rest_decoder$decode_child_imm_val$002     = decode_child_imm_val$003;
  assign rest_decoder$decode_child_op_class$000    = decode_child_op_class$001;
  assign rest_decoder$decode_child_op_class$001    = decode_child_op_class$002;
  assign rest_decoder$decode_child_op_class$002    = decode_child_op_class$003;
  assign rest_decoder$decode_child_rd_val$000      = decode_child_rd_val$001;
  assign rest_decoder$decode_child_rd_val$001      = decode_child_rd_val$002;
  assign rest_decoder$decode_child_rd_val$002      = decode_child_rd_val$003;
  assign rest_decoder$decode_child_result$000      = decode_child_result$001;
  assign rest_decoder$decode_child_result$001      = decode_child_result$002;
  assign rest_decoder$decode_child_result$002      = decode_child_result$003;
  assign rest_decoder$decode_child_rs1_val$000     = decode_child_rs1_val$001;
  assign rest_decoder$decode_child_rs1_val$001     = decode_child_rs1_val$002;
  assign rest_decoder$decode_child_rs1_val$002     = decode_child_rs1_val$003;
  assign rest_decoder$decode_child_rs2_val$000     = decode_child_rs2_val$001;
  assign rest_decoder$decode_child_rs2_val$001     = decode_child_rs2_val$002;
  assign rest_decoder$decode_child_rs2_val$002     = decode_child_rs2_val$003;
  assign rest_decoder$decode_child_serialize$000   = decode_child_serialize$001;
  assign rest_decoder$decode_child_serialize$001   = decode_child_serialize$002;
  assign rest_decoder$decode_child_serialize$002   = decode_child_serialize$003;
  assign rest_decoder$decode_child_speculative$000 = decode_child_speculative$001;
  assign rest_decoder$decode_child_speculative$001 = decode_child_speculative$002;
  assign rest_decoder$decode_child_speculative$002 = decode_child_speculative$003;
  assign rest_decoder$decode_child_success$000     = decode_child_success$001;
  assign rest_decoder$decode_child_success$001     = decode_child_success$002;
  assign rest_decoder$decode_child_success$002     = decode_child_success$003;
  assign rest_decoder$decode_inst                  = binary_decoder$decode_b_inst;
  assign rest_decoder$reset                        = reset;



endmodule // CompositeDecoder_0x2c27817f253ceafb

//-----------------------------------------------------------------------------
// CompositeDecoder_0x2c27817f250f23b4
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"nchildren": 3}
// PyMTL: verilator_xinit = zeros
module CompositeDecoder_0x2c27817f250f23b4
(
  input  logic [   0:0] clk,
  input  logic [   2:0] decode_child_imm_type$000,
  input  logic [   2:0] decode_child_imm_type$001,
  input  logic [   2:0] decode_child_imm_type$002,
  input  logic [   0:0] decode_child_imm_val$000,
  input  logic [   0:0] decode_child_imm_val$001,
  input  logic [   0:0] decode_child_imm_val$002,
  output logic [  31:0] decode_child_inst$000,
  output logic [  31:0] decode_child_inst$001,
  output logic [  31:0] decode_child_inst$002,
  input  logic [   2:0] decode_child_op_class$000,
  input  logic [   2:0] decode_child_op_class$001,
  input  logic [   2:0] decode_child_op_class$002,
  input  logic [   0:0] decode_child_rd_val$000,
  input  logic [   0:0] decode_child_rd_val$001,
  input  logic [   0:0] decode_child_rd_val$002,
  input  logic [  14:0] decode_child_result$000,
  input  logic [  14:0] decode_child_result$001,
  input  logic [  14:0] decode_child_result$002,
  input  logic [   0:0] decode_child_rs1_val$000,
  input  logic [   0:0] decode_child_rs1_val$001,
  input  logic [   0:0] decode_child_rs1_val$002,
  input  logic [   0:0] decode_child_rs2_val$000,
  input  logic [   0:0] decode_child_rs2_val$001,
  input  logic [   0:0] decode_child_rs2_val$002,
  input  logic [   0:0] decode_child_serialize$000,
  input  logic [   0:0] decode_child_serialize$001,
  input  logic [   0:0] decode_child_serialize$002,
  input  logic [   0:0] decode_child_speculative$000,
  input  logic [   0:0] decode_child_speculative$001,
  input  logic [   0:0] decode_child_speculative$002,
  input  logic [   0:0] decode_child_success$000,
  input  logic [   0:0] decode_child_success$001,
  input  logic [   0:0] decode_child_success$002,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // rest_decoder temporaries
  logic   [   0:0] rest_decoder$decode_child_serialize$000;
  logic   [   0:0] rest_decoder$decode_child_serialize$001;
  logic   [  14:0] rest_decoder$decode_child_result$000;
  logic   [  14:0] rest_decoder$decode_child_result$001;
  logic   [   0:0] rest_decoder$decode_child_imm_val$000;
  logic   [   0:0] rest_decoder$decode_child_imm_val$001;
  logic   [   0:0] rest_decoder$clk;
  logic   [   2:0] rest_decoder$decode_child_op_class$000;
  logic   [   2:0] rest_decoder$decode_child_op_class$001;
  logic   [  31:0] rest_decoder$decode_inst;
  logic   [   0:0] rest_decoder$decode_child_rd_val$000;
  logic   [   0:0] rest_decoder$decode_child_rd_val$001;
  logic   [   0:0] rest_decoder$decode_child_speculative$000;
  logic   [   0:0] rest_decoder$decode_child_speculative$001;
  logic   [   0:0] rest_decoder$decode_child_success$000;
  logic   [   0:0] rest_decoder$decode_child_success$001;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$000;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$001;
  logic   [   0:0] rest_decoder$reset;
  logic   [   2:0] rest_decoder$decode_child_imm_type$000;
  logic   [   2:0] rest_decoder$decode_child_imm_type$001;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$000;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$001;
  logic   [   2:0] rest_decoder$decode_imm_type;
  logic   [  31:0] rest_decoder$decode_child_inst$000;
  logic   [  31:0] rest_decoder$decode_child_inst$001;
  logic   [   0:0] rest_decoder$decode_serialize;
  logic   [  14:0] rest_decoder$decode_result;
  logic   [   0:0] rest_decoder$decode_imm_val;
  logic   [   0:0] rest_decoder$decode_rd_val;
  logic   [   0:0] rest_decoder$decode_rs2_val;
  logic   [   2:0] rest_decoder$decode_op_class;
  logic   [   0:0] rest_decoder$decode_success;
  logic   [   0:0] rest_decoder$decode_speculative;
  logic   [   0:0] rest_decoder$decode_rs1_val;

  CompositeDecoder_0x2c27817f251e6671 rest_decoder
  (
    .decode_child_serialize$000   ( rest_decoder$decode_child_serialize$000 ),
    .decode_child_serialize$001   ( rest_decoder$decode_child_serialize$001 ),
    .decode_child_result$000      ( rest_decoder$decode_child_result$000 ),
    .decode_child_result$001      ( rest_decoder$decode_child_result$001 ),
    .decode_child_imm_val$000     ( rest_decoder$decode_child_imm_val$000 ),
    .decode_child_imm_val$001     ( rest_decoder$decode_child_imm_val$001 ),
    .clk                          ( rest_decoder$clk ),
    .decode_child_op_class$000    ( rest_decoder$decode_child_op_class$000 ),
    .decode_child_op_class$001    ( rest_decoder$decode_child_op_class$001 ),
    .decode_inst                  ( rest_decoder$decode_inst ),
    .decode_child_rd_val$000      ( rest_decoder$decode_child_rd_val$000 ),
    .decode_child_rd_val$001      ( rest_decoder$decode_child_rd_val$001 ),
    .decode_child_speculative$000 ( rest_decoder$decode_child_speculative$000 ),
    .decode_child_speculative$001 ( rest_decoder$decode_child_speculative$001 ),
    .decode_child_success$000     ( rest_decoder$decode_child_success$000 ),
    .decode_child_success$001     ( rest_decoder$decode_child_success$001 ),
    .decode_child_rs2_val$000     ( rest_decoder$decode_child_rs2_val$000 ),
    .decode_child_rs2_val$001     ( rest_decoder$decode_child_rs2_val$001 ),
    .reset                        ( rest_decoder$reset ),
    .decode_child_imm_type$000    ( rest_decoder$decode_child_imm_type$000 ),
    .decode_child_imm_type$001    ( rest_decoder$decode_child_imm_type$001 ),
    .decode_child_rs1_val$000     ( rest_decoder$decode_child_rs1_val$000 ),
    .decode_child_rs1_val$001     ( rest_decoder$decode_child_rs1_val$001 ),
    .decode_imm_type              ( rest_decoder$decode_imm_type ),
    .decode_child_inst$000        ( rest_decoder$decode_child_inst$000 ),
    .decode_child_inst$001        ( rest_decoder$decode_child_inst$001 ),
    .decode_serialize             ( rest_decoder$decode_serialize ),
    .decode_result                ( rest_decoder$decode_result ),
    .decode_imm_val               ( rest_decoder$decode_imm_val ),
    .decode_rd_val                ( rest_decoder$decode_rd_val ),
    .decode_rs2_val               ( rest_decoder$decode_rs2_val ),
    .decode_op_class              ( rest_decoder$decode_op_class ),
    .decode_success               ( rest_decoder$decode_success ),
    .decode_speculative           ( rest_decoder$decode_speculative ),
    .decode_rs1_val               ( rest_decoder$decode_rs1_val )
  );

  // binary_decoder temporaries
  logic   [   0:0] binary_decoder$decode_b_rs1_val;
  logic   [   0:0] binary_decoder$decode_a_rs1_val;
  logic   [   0:0] binary_decoder$decode_b_rs2_val;
  logic   [   0:0] binary_decoder$decode_a_serialize;
  logic   [  14:0] binary_decoder$decode_a_result;
  logic   [   0:0] binary_decoder$clk;
  logic   [   2:0] binary_decoder$decode_a_imm_type;
  logic   [  31:0] binary_decoder$decode_inst;
  logic   [   0:0] binary_decoder$decode_b_rd_val;
  logic   [   0:0] binary_decoder$decode_a_speculative;
  logic   [   0:0] binary_decoder$decode_a_imm_val;
  logic   [   0:0] binary_decoder$decode_b_success;
  logic   [   2:0] binary_decoder$decode_a_op_class;
  logic   [   0:0] binary_decoder$reset;
  logic   [   2:0] binary_decoder$decode_b_op_class;
  logic   [   2:0] binary_decoder$decode_b_imm_type;
  logic   [   0:0] binary_decoder$decode_a_rd_val;
  logic   [   0:0] binary_decoder$decode_a_success;
  logic   [   0:0] binary_decoder$decode_b_serialize;
  logic   [   0:0] binary_decoder$decode_b_speculative;
  logic   [  14:0] binary_decoder$decode_b_result;
  logic   [   0:0] binary_decoder$decode_a_rs2_val;
  logic   [   0:0] binary_decoder$decode_b_imm_val;
  logic   [   2:0] binary_decoder$decode_imm_type;
  logic   [  31:0] binary_decoder$decode_a_inst;
  logic   [   0:0] binary_decoder$decode_serialize;
  logic   [  14:0] binary_decoder$decode_result;
  logic   [   0:0] binary_decoder$decode_imm_val;
  logic   [   0:0] binary_decoder$decode_rd_val;
  logic   [   0:0] binary_decoder$decode_rs2_val;
  logic   [   2:0] binary_decoder$decode_op_class;
  logic   [   0:0] binary_decoder$decode_success;
  logic   [   0:0] binary_decoder$decode_speculative;
  logic   [  31:0] binary_decoder$decode_b_inst;
  logic   [   0:0] binary_decoder$decode_rs1_val;

  BinaryCompositeDecoder_0x6047cbf454b06e40 binary_decoder
  (
    .decode_b_rs1_val     ( binary_decoder$decode_b_rs1_val ),
    .decode_a_rs1_val     ( binary_decoder$decode_a_rs1_val ),
    .decode_b_rs2_val     ( binary_decoder$decode_b_rs2_val ),
    .decode_a_serialize   ( binary_decoder$decode_a_serialize ),
    .decode_a_result      ( binary_decoder$decode_a_result ),
    .clk                  ( binary_decoder$clk ),
    .decode_a_imm_type    ( binary_decoder$decode_a_imm_type ),
    .decode_inst          ( binary_decoder$decode_inst ),
    .decode_b_rd_val      ( binary_decoder$decode_b_rd_val ),
    .decode_a_speculative ( binary_decoder$decode_a_speculative ),
    .decode_a_imm_val     ( binary_decoder$decode_a_imm_val ),
    .decode_b_success     ( binary_decoder$decode_b_success ),
    .decode_a_op_class    ( binary_decoder$decode_a_op_class ),
    .reset                ( binary_decoder$reset ),
    .decode_b_op_class    ( binary_decoder$decode_b_op_class ),
    .decode_b_imm_type    ( binary_decoder$decode_b_imm_type ),
    .decode_a_rd_val      ( binary_decoder$decode_a_rd_val ),
    .decode_a_success     ( binary_decoder$decode_a_success ),
    .decode_b_serialize   ( binary_decoder$decode_b_serialize ),
    .decode_b_speculative ( binary_decoder$decode_b_speculative ),
    .decode_b_result      ( binary_decoder$decode_b_result ),
    .decode_a_rs2_val     ( binary_decoder$decode_a_rs2_val ),
    .decode_b_imm_val     ( binary_decoder$decode_b_imm_val ),
    .decode_imm_type      ( binary_decoder$decode_imm_type ),
    .decode_a_inst        ( binary_decoder$decode_a_inst ),
    .decode_serialize     ( binary_decoder$decode_serialize ),
    .decode_result        ( binary_decoder$decode_result ),
    .decode_imm_val       ( binary_decoder$decode_imm_val ),
    .decode_rd_val        ( binary_decoder$decode_rd_val ),
    .decode_rs2_val       ( binary_decoder$decode_rs2_val ),
    .decode_op_class      ( binary_decoder$decode_op_class ),
    .decode_success       ( binary_decoder$decode_success ),
    .decode_speculative   ( binary_decoder$decode_speculative ),
    .decode_b_inst        ( binary_decoder$decode_b_inst ),
    .decode_rs1_val       ( binary_decoder$decode_rs1_val )
  );

  // signal connections
  assign binary_decoder$clk                        = clk;
  assign binary_decoder$decode_a_imm_type          = decode_child_imm_type$000;
  assign binary_decoder$decode_a_imm_val           = decode_child_imm_val$000;
  assign binary_decoder$decode_a_op_class          = decode_child_op_class$000;
  assign binary_decoder$decode_a_rd_val            = decode_child_rd_val$000;
  assign binary_decoder$decode_a_result            = decode_child_result$000;
  assign binary_decoder$decode_a_rs1_val           = decode_child_rs1_val$000;
  assign binary_decoder$decode_a_rs2_val           = decode_child_rs2_val$000;
  assign binary_decoder$decode_a_serialize         = decode_child_serialize$000;
  assign binary_decoder$decode_a_speculative       = decode_child_speculative$000;
  assign binary_decoder$decode_a_success           = decode_child_success$000;
  assign binary_decoder$decode_b_imm_type          = rest_decoder$decode_imm_type;
  assign binary_decoder$decode_b_imm_val           = rest_decoder$decode_imm_val;
  assign binary_decoder$decode_b_op_class          = rest_decoder$decode_op_class;
  assign binary_decoder$decode_b_rd_val            = rest_decoder$decode_rd_val;
  assign binary_decoder$decode_b_result            = rest_decoder$decode_result;
  assign binary_decoder$decode_b_rs1_val           = rest_decoder$decode_rs1_val;
  assign binary_decoder$decode_b_rs2_val           = rest_decoder$decode_rs2_val;
  assign binary_decoder$decode_b_serialize         = rest_decoder$decode_serialize;
  assign binary_decoder$decode_b_speculative       = rest_decoder$decode_speculative;
  assign binary_decoder$decode_b_success           = rest_decoder$decode_success;
  assign binary_decoder$decode_inst                = decode_inst;
  assign binary_decoder$reset                      = reset;
  assign decode_child_inst$000                     = binary_decoder$decode_a_inst;
  assign decode_child_inst$001                     = rest_decoder$decode_child_inst$000;
  assign decode_child_inst$002                     = rest_decoder$decode_child_inst$001;
  assign decode_imm_type                           = binary_decoder$decode_imm_type;
  assign decode_imm_val                            = binary_decoder$decode_imm_val;
  assign decode_op_class                           = binary_decoder$decode_op_class;
  assign decode_rd_val                             = binary_decoder$decode_rd_val;
  assign decode_result                             = binary_decoder$decode_result;
  assign decode_rs1_val                            = binary_decoder$decode_rs1_val;
  assign decode_rs2_val                            = binary_decoder$decode_rs2_val;
  assign decode_serialize                          = binary_decoder$decode_serialize;
  assign decode_speculative                        = binary_decoder$decode_speculative;
  assign decode_success                            = binary_decoder$decode_success;
  assign rest_decoder$clk                          = clk;
  assign rest_decoder$decode_child_imm_type$000    = decode_child_imm_type$001;
  assign rest_decoder$decode_child_imm_type$001    = decode_child_imm_type$002;
  assign rest_decoder$decode_child_imm_val$000     = decode_child_imm_val$001;
  assign rest_decoder$decode_child_imm_val$001     = decode_child_imm_val$002;
  assign rest_decoder$decode_child_op_class$000    = decode_child_op_class$001;
  assign rest_decoder$decode_child_op_class$001    = decode_child_op_class$002;
  assign rest_decoder$decode_child_rd_val$000      = decode_child_rd_val$001;
  assign rest_decoder$decode_child_rd_val$001      = decode_child_rd_val$002;
  assign rest_decoder$decode_child_result$000      = decode_child_result$001;
  assign rest_decoder$decode_child_result$001      = decode_child_result$002;
  assign rest_decoder$decode_child_rs1_val$000     = decode_child_rs1_val$001;
  assign rest_decoder$decode_child_rs1_val$001     = decode_child_rs1_val$002;
  assign rest_decoder$decode_child_rs2_val$000     = decode_child_rs2_val$001;
  assign rest_decoder$decode_child_rs2_val$001     = decode_child_rs2_val$002;
  assign rest_decoder$decode_child_serialize$000   = decode_child_serialize$001;
  assign rest_decoder$decode_child_serialize$001   = decode_child_serialize$002;
  assign rest_decoder$decode_child_speculative$000 = decode_child_speculative$001;
  assign rest_decoder$decode_child_speculative$001 = decode_child_speculative$002;
  assign rest_decoder$decode_child_success$000     = decode_child_success$001;
  assign rest_decoder$decode_child_success$001     = decode_child_success$002;
  assign rest_decoder$decode_inst                  = binary_decoder$decode_b_inst;
  assign rest_decoder$reset                        = reset;



endmodule // CompositeDecoder_0x2c27817f250f23b4

//-----------------------------------------------------------------------------
// CompositeDecoder_0x2c27817f251e6671
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"nchildren": 2}
// PyMTL: verilator_xinit = zeros
module CompositeDecoder_0x2c27817f251e6671
(
  input  logic [   0:0] clk,
  input  logic [   2:0] decode_child_imm_type$000,
  input  logic [   2:0] decode_child_imm_type$001,
  input  logic [   0:0] decode_child_imm_val$000,
  input  logic [   0:0] decode_child_imm_val$001,
  output logic [  31:0] decode_child_inst$000,
  output logic [  31:0] decode_child_inst$001,
  input  logic [   2:0] decode_child_op_class$000,
  input  logic [   2:0] decode_child_op_class$001,
  input  logic [   0:0] decode_child_rd_val$000,
  input  logic [   0:0] decode_child_rd_val$001,
  input  logic [  14:0] decode_child_result$000,
  input  logic [  14:0] decode_child_result$001,
  input  logic [   0:0] decode_child_rs1_val$000,
  input  logic [   0:0] decode_child_rs1_val$001,
  input  logic [   0:0] decode_child_rs2_val$000,
  input  logic [   0:0] decode_child_rs2_val$001,
  input  logic [   0:0] decode_child_serialize$000,
  input  logic [   0:0] decode_child_serialize$001,
  input  logic [   0:0] decode_child_speculative$000,
  input  logic [   0:0] decode_child_speculative$001,
  input  logic [   0:0] decode_child_success$000,
  input  logic [   0:0] decode_child_success$001,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // rest_decoder temporaries
  logic   [   0:0] rest_decoder$decode_child_serialize$000;
  logic   [  14:0] rest_decoder$decode_child_result$000;
  logic   [   0:0] rest_decoder$decode_child_imm_val$000;
  logic   [   0:0] rest_decoder$clk;
  logic   [   2:0] rest_decoder$decode_child_op_class$000;
  logic   [  31:0] rest_decoder$decode_inst;
  logic   [   0:0] rest_decoder$decode_child_rd_val$000;
  logic   [   0:0] rest_decoder$decode_child_speculative$000;
  logic   [   0:0] rest_decoder$decode_child_success$000;
  logic   [   0:0] rest_decoder$decode_child_rs2_val$000;
  logic   [   0:0] rest_decoder$reset;
  logic   [   2:0] rest_decoder$decode_child_imm_type$000;
  logic   [   0:0] rest_decoder$decode_child_rs1_val$000;
  logic   [   2:0] rest_decoder$decode_imm_type;
  logic   [  31:0] rest_decoder$decode_child_inst$000;
  logic   [   0:0] rest_decoder$decode_serialize;
  logic   [  14:0] rest_decoder$decode_result;
  logic   [   0:0] rest_decoder$decode_imm_val;
  logic   [   0:0] rest_decoder$decode_rd_val;
  logic   [   0:0] rest_decoder$decode_rs2_val;
  logic   [   2:0] rest_decoder$decode_op_class;
  logic   [   0:0] rest_decoder$decode_success;
  logic   [   0:0] rest_decoder$decode_speculative;
  logic   [   0:0] rest_decoder$decode_rs1_val;

  CompositeDecoder_0x2c27817f24f09f0a rest_decoder
  (
    .decode_child_serialize$000   ( rest_decoder$decode_child_serialize$000 ),
    .decode_child_result$000      ( rest_decoder$decode_child_result$000 ),
    .decode_child_imm_val$000     ( rest_decoder$decode_child_imm_val$000 ),
    .clk                          ( rest_decoder$clk ),
    .decode_child_op_class$000    ( rest_decoder$decode_child_op_class$000 ),
    .decode_inst                  ( rest_decoder$decode_inst ),
    .decode_child_rd_val$000      ( rest_decoder$decode_child_rd_val$000 ),
    .decode_child_speculative$000 ( rest_decoder$decode_child_speculative$000 ),
    .decode_child_success$000     ( rest_decoder$decode_child_success$000 ),
    .decode_child_rs2_val$000     ( rest_decoder$decode_child_rs2_val$000 ),
    .reset                        ( rest_decoder$reset ),
    .decode_child_imm_type$000    ( rest_decoder$decode_child_imm_type$000 ),
    .decode_child_rs1_val$000     ( rest_decoder$decode_child_rs1_val$000 ),
    .decode_imm_type              ( rest_decoder$decode_imm_type ),
    .decode_child_inst$000        ( rest_decoder$decode_child_inst$000 ),
    .decode_serialize             ( rest_decoder$decode_serialize ),
    .decode_result                ( rest_decoder$decode_result ),
    .decode_imm_val               ( rest_decoder$decode_imm_val ),
    .decode_rd_val                ( rest_decoder$decode_rd_val ),
    .decode_rs2_val               ( rest_decoder$decode_rs2_val ),
    .decode_op_class              ( rest_decoder$decode_op_class ),
    .decode_success               ( rest_decoder$decode_success ),
    .decode_speculative           ( rest_decoder$decode_speculative ),
    .decode_rs1_val               ( rest_decoder$decode_rs1_val )
  );

  // binary_decoder temporaries
  logic   [   0:0] binary_decoder$decode_b_rs1_val;
  logic   [   0:0] binary_decoder$decode_a_rs1_val;
  logic   [   0:0] binary_decoder$decode_b_rs2_val;
  logic   [   0:0] binary_decoder$decode_a_serialize;
  logic   [  14:0] binary_decoder$decode_a_result;
  logic   [   0:0] binary_decoder$clk;
  logic   [   2:0] binary_decoder$decode_a_imm_type;
  logic   [  31:0] binary_decoder$decode_inst;
  logic   [   0:0] binary_decoder$decode_b_rd_val;
  logic   [   0:0] binary_decoder$decode_a_speculative;
  logic   [   0:0] binary_decoder$decode_a_imm_val;
  logic   [   0:0] binary_decoder$decode_b_success;
  logic   [   2:0] binary_decoder$decode_a_op_class;
  logic   [   0:0] binary_decoder$reset;
  logic   [   2:0] binary_decoder$decode_b_op_class;
  logic   [   2:0] binary_decoder$decode_b_imm_type;
  logic   [   0:0] binary_decoder$decode_a_rd_val;
  logic   [   0:0] binary_decoder$decode_a_success;
  logic   [   0:0] binary_decoder$decode_b_serialize;
  logic   [   0:0] binary_decoder$decode_b_speculative;
  logic   [  14:0] binary_decoder$decode_b_result;
  logic   [   0:0] binary_decoder$decode_a_rs2_val;
  logic   [   0:0] binary_decoder$decode_b_imm_val;
  logic   [   2:0] binary_decoder$decode_imm_type;
  logic   [  31:0] binary_decoder$decode_a_inst;
  logic   [   0:0] binary_decoder$decode_serialize;
  logic   [  14:0] binary_decoder$decode_result;
  logic   [   0:0] binary_decoder$decode_imm_val;
  logic   [   0:0] binary_decoder$decode_rd_val;
  logic   [   0:0] binary_decoder$decode_rs2_val;
  logic   [   2:0] binary_decoder$decode_op_class;
  logic   [   0:0] binary_decoder$decode_success;
  logic   [   0:0] binary_decoder$decode_speculative;
  logic   [  31:0] binary_decoder$decode_b_inst;
  logic   [   0:0] binary_decoder$decode_rs1_val;

  BinaryCompositeDecoder_0x6047cbf454b06e40 binary_decoder
  (
    .decode_b_rs1_val     ( binary_decoder$decode_b_rs1_val ),
    .decode_a_rs1_val     ( binary_decoder$decode_a_rs1_val ),
    .decode_b_rs2_val     ( binary_decoder$decode_b_rs2_val ),
    .decode_a_serialize   ( binary_decoder$decode_a_serialize ),
    .decode_a_result      ( binary_decoder$decode_a_result ),
    .clk                  ( binary_decoder$clk ),
    .decode_a_imm_type    ( binary_decoder$decode_a_imm_type ),
    .decode_inst          ( binary_decoder$decode_inst ),
    .decode_b_rd_val      ( binary_decoder$decode_b_rd_val ),
    .decode_a_speculative ( binary_decoder$decode_a_speculative ),
    .decode_a_imm_val     ( binary_decoder$decode_a_imm_val ),
    .decode_b_success     ( binary_decoder$decode_b_success ),
    .decode_a_op_class    ( binary_decoder$decode_a_op_class ),
    .reset                ( binary_decoder$reset ),
    .decode_b_op_class    ( binary_decoder$decode_b_op_class ),
    .decode_b_imm_type    ( binary_decoder$decode_b_imm_type ),
    .decode_a_rd_val      ( binary_decoder$decode_a_rd_val ),
    .decode_a_success     ( binary_decoder$decode_a_success ),
    .decode_b_serialize   ( binary_decoder$decode_b_serialize ),
    .decode_b_speculative ( binary_decoder$decode_b_speculative ),
    .decode_b_result      ( binary_decoder$decode_b_result ),
    .decode_a_rs2_val     ( binary_decoder$decode_a_rs2_val ),
    .decode_b_imm_val     ( binary_decoder$decode_b_imm_val ),
    .decode_imm_type      ( binary_decoder$decode_imm_type ),
    .decode_a_inst        ( binary_decoder$decode_a_inst ),
    .decode_serialize     ( binary_decoder$decode_serialize ),
    .decode_result        ( binary_decoder$decode_result ),
    .decode_imm_val       ( binary_decoder$decode_imm_val ),
    .decode_rd_val        ( binary_decoder$decode_rd_val ),
    .decode_rs2_val       ( binary_decoder$decode_rs2_val ),
    .decode_op_class      ( binary_decoder$decode_op_class ),
    .decode_success       ( binary_decoder$decode_success ),
    .decode_speculative   ( binary_decoder$decode_speculative ),
    .decode_b_inst        ( binary_decoder$decode_b_inst ),
    .decode_rs1_val       ( binary_decoder$decode_rs1_val )
  );

  // signal connections
  assign binary_decoder$clk                        = clk;
  assign binary_decoder$decode_a_imm_type          = decode_child_imm_type$000;
  assign binary_decoder$decode_a_imm_val           = decode_child_imm_val$000;
  assign binary_decoder$decode_a_op_class          = decode_child_op_class$000;
  assign binary_decoder$decode_a_rd_val            = decode_child_rd_val$000;
  assign binary_decoder$decode_a_result            = decode_child_result$000;
  assign binary_decoder$decode_a_rs1_val           = decode_child_rs1_val$000;
  assign binary_decoder$decode_a_rs2_val           = decode_child_rs2_val$000;
  assign binary_decoder$decode_a_serialize         = decode_child_serialize$000;
  assign binary_decoder$decode_a_speculative       = decode_child_speculative$000;
  assign binary_decoder$decode_a_success           = decode_child_success$000;
  assign binary_decoder$decode_b_imm_type          = rest_decoder$decode_imm_type;
  assign binary_decoder$decode_b_imm_val           = rest_decoder$decode_imm_val;
  assign binary_decoder$decode_b_op_class          = rest_decoder$decode_op_class;
  assign binary_decoder$decode_b_rd_val            = rest_decoder$decode_rd_val;
  assign binary_decoder$decode_b_result            = rest_decoder$decode_result;
  assign binary_decoder$decode_b_rs1_val           = rest_decoder$decode_rs1_val;
  assign binary_decoder$decode_b_rs2_val           = rest_decoder$decode_rs2_val;
  assign binary_decoder$decode_b_serialize         = rest_decoder$decode_serialize;
  assign binary_decoder$decode_b_speculative       = rest_decoder$decode_speculative;
  assign binary_decoder$decode_b_success           = rest_decoder$decode_success;
  assign binary_decoder$decode_inst                = decode_inst;
  assign binary_decoder$reset                      = reset;
  assign decode_child_inst$000                     = binary_decoder$decode_a_inst;
  assign decode_child_inst$001                     = rest_decoder$decode_child_inst$000;
  assign decode_imm_type                           = binary_decoder$decode_imm_type;
  assign decode_imm_val                            = binary_decoder$decode_imm_val;
  assign decode_op_class                           = binary_decoder$decode_op_class;
  assign decode_rd_val                             = binary_decoder$decode_rd_val;
  assign decode_result                             = binary_decoder$decode_result;
  assign decode_rs1_val                            = binary_decoder$decode_rs1_val;
  assign decode_rs2_val                            = binary_decoder$decode_rs2_val;
  assign decode_serialize                          = binary_decoder$decode_serialize;
  assign decode_speculative                        = binary_decoder$decode_speculative;
  assign decode_success                            = binary_decoder$decode_success;
  assign rest_decoder$clk                          = clk;
  assign rest_decoder$decode_child_imm_type$000    = decode_child_imm_type$001;
  assign rest_decoder$decode_child_imm_val$000     = decode_child_imm_val$001;
  assign rest_decoder$decode_child_op_class$000    = decode_child_op_class$001;
  assign rest_decoder$decode_child_rd_val$000      = decode_child_rd_val$001;
  assign rest_decoder$decode_child_result$000      = decode_child_result$001;
  assign rest_decoder$decode_child_rs1_val$000     = decode_child_rs1_val$001;
  assign rest_decoder$decode_child_rs2_val$000     = decode_child_rs2_val$001;
  assign rest_decoder$decode_child_serialize$000   = decode_child_serialize$001;
  assign rest_decoder$decode_child_speculative$000 = decode_child_speculative$001;
  assign rest_decoder$decode_child_success$000     = decode_child_success$001;
  assign rest_decoder$decode_inst                  = binary_decoder$decode_b_inst;
  assign rest_decoder$reset                        = reset;



endmodule // CompositeDecoder_0x2c27817f251e6671

//-----------------------------------------------------------------------------
// CompositeDecoder_0x2c27817f24f09f0a
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"nchildren": 1}
// PyMTL: verilator_xinit = zeros
module CompositeDecoder_0x2c27817f24f09f0a
(
  input  logic [   0:0] clk,
  input  logic [   2:0] decode_child_imm_type$000,
  input  logic [   0:0] decode_child_imm_val$000,
  output logic [  31:0] decode_child_inst$000,
  input  logic [   2:0] decode_child_op_class$000,
  input  logic [   0:0] decode_child_rd_val$000,
  input  logic [  14:0] decode_child_result$000,
  input  logic [   0:0] decode_child_rs1_val$000,
  input  logic [   0:0] decode_child_rs2_val$000,
  input  logic [   0:0] decode_child_serialize$000,
  input  logic [   0:0] decode_child_speculative$000,
  input  logic [   0:0] decode_child_success$000,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // signal connections
  assign decode_child_inst$000 = decode_inst;
  assign decode_imm_type       = decode_child_imm_type$000;
  assign decode_imm_val        = decode_child_imm_val$000;
  assign decode_op_class       = decode_child_op_class$000;
  assign decode_rd_val         = decode_child_rd_val$000;
  assign decode_result         = decode_child_result$000;
  assign decode_rs1_val        = decode_child_rs1_val$000;
  assign decode_rs2_val        = decode_child_rs2_val$000;
  assign decode_serialize      = decode_child_serialize$000;
  assign decode_speculative    = decode_child_speculative$000;
  assign decode_success        = decode_child_success$000;



endmodule // CompositeDecoder_0x2c27817f24f09f0a

//-----------------------------------------------------------------------------
// BinaryCompositeDecoder_0x6047cbf454b06e40
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {}
// PyMTL: verilator_xinit = zeros
module BinaryCompositeDecoder_0x6047cbf454b06e40
(
  input  logic [   0:0] clk,
  input  logic [   2:0] decode_a_imm_type,
  input  logic [   0:0] decode_a_imm_val,
  output logic [  31:0] decode_a_inst,
  input  logic [   2:0] decode_a_op_class,
  input  logic [   0:0] decode_a_rd_val,
  input  logic [  14:0] decode_a_result,
  input  logic [   0:0] decode_a_rs1_val,
  input  logic [   0:0] decode_a_rs2_val,
  input  logic [   0:0] decode_a_serialize,
  input  logic [   0:0] decode_a_speculative,
  input  logic [   0:0] decode_a_success,
  input  logic [   2:0] decode_b_imm_type,
  input  logic [   0:0] decode_b_imm_val,
  output logic [  31:0] decode_b_inst,
  input  logic [   2:0] decode_b_op_class,
  input  logic [   0:0] decode_b_rd_val,
  input  logic [  14:0] decode_b_result,
  input  logic [   0:0] decode_b_rs1_val,
  input  logic [   0:0] decode_b_rs2_val,
  input  logic [   0:0] decode_b_serialize,
  input  logic [   0:0] decode_b_speculative,
  input  logic [   0:0] decode_b_success,
  output logic  [   2:0] decode_imm_type,
  output logic  [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic  [   2:0] decode_op_class,
  output logic  [   0:0] decode_rd_val,
  output logic  [  14:0] decode_result,
  output logic  [   0:0] decode_rs1_val,
  output logic  [   0:0] decode_rs2_val,
  output logic  [   0:0] decode_serialize,
  output logic  [   0:0] decode_speculative,
  output logic  [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // signal connections
  assign decode_a_inst = decode_inst;
  assign decode_b_inst = decode_inst;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pick():
  //       if s.decode_a_success:
  //         s.decode_success.v = s.decode_a_success
  //         s.decode_serialize.v = s.decode_a_serialize
  //         s.decode_speculative.v = s.decode_a_speculative
  //         s.decode_rs1_val.v = s.decode_a_rs1_val
  //         s.decode_rs2_val.v = s.decode_a_rs2_val
  //         s.decode_rd_val.v = s.decode_a_rd_val
  //         s.decode_imm_type.v = s.decode_a_imm_type
  //         s.decode_imm_val.v = s.decode_a_imm_val
  //         s.decode_op_class.v = s.decode_a_op_class
  //         s.decode_result.v = s.decode_a_result
  //       else:
  //         s.decode_success.v = s.decode_b_success
  //         s.decode_serialize.v = s.decode_b_serialize
  //         s.decode_speculative.v = s.decode_b_speculative
  //         s.decode_rs1_val.v = s.decode_b_rs1_val
  //         s.decode_rs2_val.v = s.decode_b_rs2_val
  //         s.decode_rd_val.v = s.decode_b_rd_val
  //         s.decode_imm_type.v = s.decode_b_imm_type
  //         s.decode_imm_val.v = s.decode_b_imm_val
  //         s.decode_op_class.v = s.decode_b_op_class
  //         s.decode_result.v = s.decode_b_result

  // logic for pick()
  always @ (*) begin
    if (decode_a_success) begin
      decode_success = decode_a_success;
      decode_serialize = decode_a_serialize;
      decode_speculative = decode_a_speculative;
      decode_rs1_val = decode_a_rs1_val;
      decode_rs2_val = decode_a_rs2_val;
      decode_rd_val = decode_a_rd_val;
      decode_imm_type = decode_a_imm_type;
      decode_imm_val = decode_a_imm_val;
      decode_op_class = decode_a_op_class;
      decode_result = decode_a_result;
    end
    else begin
      decode_success = decode_b_success;
      decode_serialize = decode_b_serialize;
      decode_speculative = decode_b_speculative;
      decode_rs1_val = decode_b_rs1_val;
      decode_rs2_val = decode_b_rs2_val;
      decode_rd_val = decode_b_rd_val;
      decode_imm_type = decode_b_imm_type;
      decode_imm_val = decode_b_imm_val;
      decode_op_class = decode_b_op_class;
      decode_result = decode_b_result;
    end
  end


endmodule // BinaryCompositeDecoder_0x6047cbf454b06e40

//-----------------------------------------------------------------------------
// CsrDecoder_0x39519b5cedf33556
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.csr_decoder {}
// PyMTL: verilator_xinit = zeros
module CsrDecoder_0x39519b5cedf33556
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // generator temporaries
  logic   [  31:0] generator$gen_inst;
  logic   [   1:0] generator$gen_data;
  logic   [   0:0] generator$clk;
  logic   [   0:0] generator$reset;
  logic   [  14:0] generator$gen_payload;
  logic   [   0:0] generator$gen_valid;

  CsrPayloadGenerator_0x39519b5cedf33556 generator
  (
    .gen_inst    ( generator$gen_inst ),
    .gen_data    ( generator$gen_data ),
    .clk         ( generator$clk ),
    .reset       ( generator$reset ),
    .gen_payload ( generator$gen_payload ),
    .gen_valid   ( generator$gen_valid )
  );

  // decoder temporaries
  logic   [   0:0] decoder$clk;
  logic   [  14:0] decoder$gen_payload;
  logic   [  31:0] decoder$decode_inst;
  logic   [   0:0] decoder$gen_valid;
  logic   [   0:0] decoder$reset;
  logic   [  31:0] decoder$gen_inst;
  logic   [   2:0] decoder$decode_imm_type;
  logic   [   1:0] decoder$gen_data;
  logic   [   0:0] decoder$decode_serialize;
  logic   [  14:0] decoder$decode_result;
  logic   [   0:0] decoder$decode_imm_val;
  logic   [   0:0] decoder$decode_rd_val;
  logic   [   0:0] decoder$decode_rs2_val;
  logic   [   2:0] decoder$decode_op_class;
  logic   [   0:0] decoder$decode_success;
  logic   [   0:0] decoder$decode_speculative;
  logic   [   0:0] decoder$decode_rs1_val;

  GenDecoder_0x68c1274fba277f87 decoder
  (
    .clk                ( decoder$clk ),
    .gen_payload        ( decoder$gen_payload ),
    .decode_inst        ( decoder$decode_inst ),
    .gen_valid          ( decoder$gen_valid ),
    .reset              ( decoder$reset ),
    .gen_inst           ( decoder$gen_inst ),
    .decode_imm_type    ( decoder$decode_imm_type ),
    .gen_data           ( decoder$gen_data ),
    .decode_serialize   ( decoder$decode_serialize ),
    .decode_result      ( decoder$decode_result ),
    .decode_imm_val     ( decoder$decode_imm_val ),
    .decode_rd_val      ( decoder$decode_rd_val ),
    .decode_rs2_val     ( decoder$decode_rs2_val ),
    .decode_op_class    ( decoder$decode_op_class ),
    .decode_success     ( decoder$decode_success ),
    .decode_speculative ( decoder$decode_speculative ),
    .decode_rs1_val     ( decoder$decode_rs1_val )
  );

  // signal connections
  assign decode_imm_type     = decoder$decode_imm_type;
  assign decode_imm_val      = decoder$decode_imm_val;
  assign decode_op_class     = decoder$decode_op_class;
  assign decode_rd_val       = decoder$decode_rd_val;
  assign decode_result       = decoder$decode_result;
  assign decode_rs1_val      = decoder$decode_rs1_val;
  assign decode_rs2_val      = decoder$decode_rs2_val;
  assign decode_serialize    = decoder$decode_serialize;
  assign decode_speculative  = decoder$decode_speculative;
  assign decode_success      = decoder$decode_success;
  assign decoder$clk         = clk;
  assign decoder$decode_inst = decode_inst;
  assign decoder$gen_payload = generator$gen_payload;
  assign decoder$gen_valid   = generator$gen_valid;
  assign decoder$reset       = reset;
  assign generator$clk       = clk;
  assign generator$gen_data  = decoder$gen_data;
  assign generator$gen_inst  = decoder$gen_inst;
  assign generator$reset     = reset;



endmodule // CsrDecoder_0x39519b5cedf33556

//-----------------------------------------------------------------------------
// CsrPayloadGenerator_0x39519b5cedf33556
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.csr_decoder {}
// PyMTL: verilator_xinit = zeros
module CsrPayloadGenerator_0x39519b5cedf33556
(
  input  logic [   0:0] clk,
  input  logic [   1:0] gen_data,
  input  logic [  31:0] gen_inst,
  output logic  [  14:0] gen_payload,
  output logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // signal connections
  assign gen_valid = 1'd1;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def check_rs1_is_x0():
  //       s.gen_payload.func.v = s.gen_data
  //       s.gen_payload.csr_num.v = s.gen_inst.csrnum
  //       s.gen_payload.rs1_is_x0.v = (s.gen_inst.rs1 == 0)

  // logic for check_rs1_is_x0()
  always @ (*) begin
    gen_payload[(2)-1:0] = gen_data;
    gen_payload[(14)-1:2] = gen_inst[(32)-1:20];
    gen_payload[(15)-1:14] = (gen_inst[(20)-1:15] == 0);
  end


endmodule // CsrPayloadGenerator_0x39519b5cedf33556

//-----------------------------------------------------------------------------
// GenDecoder_0x68c1274fba277f87
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"In": 2, "ResultKind": 15, "field_list": ["funct3"], "field_map": {"1": "0", "2": "1", "3": "2"}, "fixed_map": {"opcode": "73"}, "imm_type": 0, "imm_val": 0, "op_class": 3, "rd_val": 1, "result_field": "csr_msg", "rs1_val": 1, "rs2_val": 0, "serialize": 1, "speculative": 0}
// PyMTL: verilator_xinit = zeros
module GenDecoder_0x68c1274fba277f87
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic  [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic  [   0:0] decode_success,
  output logic [   1:0] gen_data,
  output logic [  31:0] gen_inst,
  input  logic [  14:0] gen_payload,
  input  logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] fixed_equals$000;
  logic   [   1:0] lookup_out;


  // lut temporaries
  logic   [   0:0] lut$clk;
  logic   [   0:0] lut$reset;
  logic   [   2:0] lut$lookup_in_;
  logic   [   1:0] lut$lookup_out;
  logic   [   0:0] lut$lookup_valid;

  LookupTable_0x65c646caf3c5c188 lut
  (
    .clk          ( lut$clk ),
    .reset        ( lut$reset ),
    .lookup_in_   ( lut$lookup_in_ ),
    .lookup_out   ( lut$lookup_out ),
    .lookup_valid ( lut$lookup_valid )
  );

  // equals_units$000 temporaries
  logic   [   0:0] equals_units$000$clk;
  logic   [   6:0] equals_units$000$compare_in_a;
  logic   [   6:0] equals_units$000$compare_in_b;
  logic   [   0:0] equals_units$000$reset;
  logic   [   0:0] equals_units$000$compare_out;

  Equals_0x6924ce1fe1e63d28 equals_units$000
  (
    .clk          ( equals_units$000$clk ),
    .compare_in_a ( equals_units$000$compare_in_a ),
    .compare_in_b ( equals_units$000$compare_in_b ),
    .reset        ( equals_units$000$reset ),
    .compare_out  ( equals_units$000$compare_out )
  );

  // and_unit temporaries
  logic   [   0:0] and_unit$op_in_$000;
  logic   [   0:0] and_unit$op_in_$001;
  logic   [   0:0] and_unit$clk;
  logic   [   0:0] and_unit$reset;
  logic   [   0:0] and_unit$op_out;

  And_0x8e49eae68bebab2 and_unit
  (
    .op_in_$000 ( and_unit$op_in_$000 ),
    .op_in_$001 ( and_unit$op_in_$001 ),
    .clk        ( and_unit$clk ),
    .reset      ( and_unit$reset ),
    .op_out     ( and_unit$op_out )
  );

  // signal connections
  assign and_unit$clk                  = clk;
  assign and_unit$op_in_$000           = equals_units$000$compare_out;
  assign and_unit$op_in_$001           = lut$lookup_valid;
  assign and_unit$reset                = reset;
  assign decode_imm_type               = 3'd0;
  assign decode_imm_val                = 1'd0;
  assign decode_op_class               = 3'd3;
  assign decode_rd_val                 = 1'd1;
  assign decode_rs1_val                = 1'd1;
  assign decode_rs2_val                = 1'd0;
  assign decode_serialize              = 1'd1;
  assign decode_speculative            = 1'd0;
  assign equals_units$000$clk          = clk;
  assign equals_units$000$compare_in_a = decode_inst[6:0];
  assign equals_units$000$compare_in_b = 7'd115;
  assign equals_units$000$reset        = reset;
  assign gen_data                      = lookup_out;
  assign gen_inst                      = decode_inst;
  assign lookup_out                    = lut$lookup_out;
  assign lut$clk                       = clk;
  assign lut$lookup_in_[2:0]           = decode_inst[14:12];
  assign lut$reset                     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_result(rs=result_field_slice.start, re=result_field_slice.stop):
  //       s.decode_result.v = 0
  //       s.decode_result[rs:re].v = s.gen_payload

  // logic for connect_result()
  always @ (*) begin
    decode_result = 0;
    decode_result[(15)-1:0] = gen_payload;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_success():
  //       s.decode_success.v = s.gen_valid & s.and_unit.op_out

  // logic for compute_success()
  always @ (*) begin
    decode_success = (gen_valid&and_unit$op_out);
  end


endmodule // GenDecoder_0x68c1274fba277f87

//-----------------------------------------------------------------------------
// LookupTable_0x65c646caf3c5c188
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(3)) -> (valid: Bits(1), out: Bits(2))", "mapping": {"1": "0", "2": "1", "3": "2"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0x65c646caf3c5c188
(
  input  logic [   0:0] clk,
  input  logic [   2:0] lookup_in_,
  output logic [   1:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   1:0] mux$mux_default;
  logic   [   1:0] mux$mux_in_$000;
  logic   [   1:0] mux$mux_in_$001;
  logic   [   1:0] mux$mux_in_$002;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   2:0] mux$mux_select;
  logic   [   1:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x664196ff7afb375b mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 2'd0;
  assign mux$mux_in_$000 = 2'd0;
  assign mux$mux_in_$001 = 2'd1;
  assign mux$mux_in_$002 = 2'd2;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0x65c646caf3c5c188

//-----------------------------------------------------------------------------
// CaseMux_0x664196ff7afb375b
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(2), in_: Bits(2) [3], select: Bits(3)) -> (out: Bits(2), matched: Bits(1))", "svalues": ["1", "2", "3"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x664196ff7afb375b
(
  input  logic [   0:0] clk,
  input  logic [   1:0] mux_default,
  input  logic [   1:0] mux_in_$000,
  input  logic [   1:0] mux_in_$001,
  input  logic [   1:0] mux_in_$002,
  output logic [   0:0] mux_matched,
  output logic [   1:0] mux_out,
  input  logic [   2:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   1:0] out_chain$000;
  logic   [   1:0] out_chain$001;
  logic   [   1:0] out_chain$002;
  logic   [   1:0] out_chain$003;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;
  logic   [   0:0] valid_chain$003;


  // signal connections
  assign mux_matched     = valid_chain$003;
  assign mux_out         = out_chain$003;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   1:0] mux_in_[0:2];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  logic    [   1:0] out_chain[0:3];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  assign out_chain$003 = out_chain[  3];
  logic    [   0:0] valid_chain[0:3];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];
  assign valid_chain$003 = valid_chain[  3];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 1)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 2)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 3)) begin
      out_chain[3] = mux_in_[2];
      valid_chain[3] = 1;
    end
    else begin
      out_chain[3] = out_chain[2];
      valid_chain[3] = valid_chain[2];
    end
  end


endmodule // CaseMux_0x664196ff7afb375b

//-----------------------------------------------------------------------------
// GenDecoderFixed_0x30e34b165e6ab78
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"ResultKind": 3, "field_list": ["funct3"], "field_map": {"0": "type_=0x0:unsigned=0x0", "1": "type_=0x1:unsigned=0x0", "4": "type_=0x2:unsigned=0x0", "5": "type_=0x3:unsigned=0x0", "6": "type_=0x2:unsigned=0x1", "7": "type_=0x3:unsigned=0x1"}, "fixed_map": {"opcode": "63"}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 0, "result_field": "branch_msg", "rs1_val": 1, "rs2_val": 1, "serialize": 0, "speculative": 1}
// PyMTL: verilator_xinit = zeros
module GenDecoderFixed_0x30e34b165e6ab78
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic [   0:0] decode_success,
  input  logic [   0:0] reset
);

  // identity_generator temporaries
  logic   [  31:0] identity_generator$gen_inst;
  logic   [   2:0] identity_generator$gen_data;
  logic   [   0:0] identity_generator$clk;
  logic   [   0:0] identity_generator$reset;
  logic   [   2:0] identity_generator$gen_payload;
  logic   [   0:0] identity_generator$gen_valid;

  IdentityPayloadGenerator_0x56c929f0f987fa52 identity_generator
  (
    .gen_inst    ( identity_generator$gen_inst ),
    .gen_data    ( identity_generator$gen_data ),
    .clk         ( identity_generator$clk ),
    .reset       ( identity_generator$reset ),
    .gen_payload ( identity_generator$gen_payload ),
    .gen_valid   ( identity_generator$gen_valid )
  );

  // decoder temporaries
  logic   [   0:0] decoder$clk;
  logic   [   2:0] decoder$gen_payload;
  logic   [  31:0] decoder$decode_inst;
  logic   [   0:0] decoder$gen_valid;
  logic   [   0:0] decoder$reset;
  logic   [  31:0] decoder$gen_inst;
  logic   [   2:0] decoder$decode_imm_type;
  logic   [   2:0] decoder$gen_data;
  logic   [   0:0] decoder$decode_serialize;
  logic   [  14:0] decoder$decode_result;
  logic   [   0:0] decoder$decode_imm_val;
  logic   [   0:0] decoder$decode_rd_val;
  logic   [   0:0] decoder$decode_rs2_val;
  logic   [   2:0] decoder$decode_op_class;
  logic   [   0:0] decoder$decode_success;
  logic   [   0:0] decoder$decode_speculative;
  logic   [   0:0] decoder$decode_rs1_val;

  GenDecoder_0x687c848ae02befc7 decoder
  (
    .clk                ( decoder$clk ),
    .gen_payload        ( decoder$gen_payload ),
    .decode_inst        ( decoder$decode_inst ),
    .gen_valid          ( decoder$gen_valid ),
    .reset              ( decoder$reset ),
    .gen_inst           ( decoder$gen_inst ),
    .decode_imm_type    ( decoder$decode_imm_type ),
    .gen_data           ( decoder$gen_data ),
    .decode_serialize   ( decoder$decode_serialize ),
    .decode_result      ( decoder$decode_result ),
    .decode_imm_val     ( decoder$decode_imm_val ),
    .decode_rd_val      ( decoder$decode_rd_val ),
    .decode_rs2_val     ( decoder$decode_rs2_val ),
    .decode_op_class    ( decoder$decode_op_class ),
    .decode_success     ( decoder$decode_success ),
    .decode_speculative ( decoder$decode_speculative ),
    .decode_rs1_val     ( decoder$decode_rs1_val )
  );

  // signal connections
  assign decode_imm_type             = decoder$decode_imm_type;
  assign decode_imm_val              = decoder$decode_imm_val;
  assign decode_op_class             = decoder$decode_op_class;
  assign decode_rd_val               = decoder$decode_rd_val;
  assign decode_result               = decoder$decode_result;
  assign decode_rs1_val              = decoder$decode_rs1_val;
  assign decode_rs2_val              = decoder$decode_rs2_val;
  assign decode_serialize            = decoder$decode_serialize;
  assign decode_speculative          = decoder$decode_speculative;
  assign decode_success              = decoder$decode_success;
  assign decoder$clk                 = clk;
  assign decoder$decode_inst         = decode_inst;
  assign decoder$gen_payload         = identity_generator$gen_payload;
  assign decoder$gen_valid           = identity_generator$gen_valid;
  assign decoder$reset               = reset;
  assign identity_generator$clk      = clk;
  assign identity_generator$gen_data = decoder$gen_data;
  assign identity_generator$gen_inst = decoder$gen_inst;
  assign identity_generator$reset    = reset;



endmodule // GenDecoderFixed_0x30e34b165e6ab78

//-----------------------------------------------------------------------------
// IdentityPayloadGenerator_0x56c929f0f987fa52
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"interface": "gen (inst: Bits(32), data: Bits(3)) -> (valid: Bits(1), payload: Bits(3))"}
// PyMTL: verilator_xinit = zeros
module IdentityPayloadGenerator_0x56c929f0f987fa52
(
  input  logic [   0:0] clk,
  input  logic [   2:0] gen_data,
  input  logic [  31:0] gen_inst,
  output logic [   2:0] gen_payload,
  output logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // signal connections
  assign gen_payload = gen_data;
  assign gen_valid   = 1'd1;



endmodule // IdentityPayloadGenerator_0x56c929f0f987fa52

//-----------------------------------------------------------------------------
// GenDecoder_0x687c848ae02befc7
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.sub_decoder {"In": 3, "ResultKind": 3, "field_list": ["funct3"], "field_map": {"0": "type_=0x0:unsigned=0x0", "1": "type_=0x1:unsigned=0x0", "4": "type_=0x2:unsigned=0x0", "5": "type_=0x3:unsigned=0x0", "6": "type_=0x2:unsigned=0x1", "7": "type_=0x3:unsigned=0x1"}, "fixed_map": {"opcode": "63"}, "imm_type": 3, "imm_val": 1, "op_class": 3, "rd_val": 0, "result_field": "branch_msg", "rs1_val": 1, "rs2_val": 1, "serialize": 0, "speculative": 1}
// PyMTL: verilator_xinit = zeros
module GenDecoder_0x687c848ae02befc7
(
  input  logic [   0:0] clk,
  output logic [   2:0] decode_imm_type,
  output logic [   0:0] decode_imm_val,
  input  logic [  31:0] decode_inst,
  output logic [   2:0] decode_op_class,
  output logic [   0:0] decode_rd_val,
  output logic  [  14:0] decode_result,
  output logic [   0:0] decode_rs1_val,
  output logic [   0:0] decode_rs2_val,
  output logic [   0:0] decode_serialize,
  output logic [   0:0] decode_speculative,
  output logic  [   0:0] decode_success,
  output logic [   2:0] gen_data,
  output logic [  31:0] gen_inst,
  input  logic [   2:0] gen_payload,
  input  logic [   0:0] gen_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] fixed_equals$000;
  logic   [   2:0] lookup_out;


  // lut temporaries
  logic   [   0:0] lut$clk;
  logic   [   0:0] lut$reset;
  logic   [   2:0] lut$lookup_in_;
  logic   [   2:0] lut$lookup_out;
  logic   [   0:0] lut$lookup_valid;

  LookupTable_0x7098a106e042a7dc lut
  (
    .clk          ( lut$clk ),
    .reset        ( lut$reset ),
    .lookup_in_   ( lut$lookup_in_ ),
    .lookup_out   ( lut$lookup_out ),
    .lookup_valid ( lut$lookup_valid )
  );

  // equals_units$000 temporaries
  logic   [   0:0] equals_units$000$clk;
  logic   [   6:0] equals_units$000$compare_in_a;
  logic   [   6:0] equals_units$000$compare_in_b;
  logic   [   0:0] equals_units$000$reset;
  logic   [   0:0] equals_units$000$compare_out;

  Equals_0x6924ce1fe1e63d28 equals_units$000
  (
    .clk          ( equals_units$000$clk ),
    .compare_in_a ( equals_units$000$compare_in_a ),
    .compare_in_b ( equals_units$000$compare_in_b ),
    .reset        ( equals_units$000$reset ),
    .compare_out  ( equals_units$000$compare_out )
  );

  // and_unit temporaries
  logic   [   0:0] and_unit$op_in_$000;
  logic   [   0:0] and_unit$op_in_$001;
  logic   [   0:0] and_unit$clk;
  logic   [   0:0] and_unit$reset;
  logic   [   0:0] and_unit$op_out;

  And_0x8e49eae68bebab2 and_unit
  (
    .op_in_$000 ( and_unit$op_in_$000 ),
    .op_in_$001 ( and_unit$op_in_$001 ),
    .clk        ( and_unit$clk ),
    .reset      ( and_unit$reset ),
    .op_out     ( and_unit$op_out )
  );

  // signal connections
  assign and_unit$clk                  = clk;
  assign and_unit$op_in_$000           = equals_units$000$compare_out;
  assign and_unit$op_in_$001           = lut$lookup_valid;
  assign and_unit$reset                = reset;
  assign decode_imm_type               = 3'd2;
  assign decode_imm_val                = 1'd1;
  assign decode_op_class               = 3'd2;
  assign decode_rd_val                 = 1'd0;
  assign decode_rs1_val                = 1'd1;
  assign decode_rs2_val                = 1'd1;
  assign decode_serialize              = 1'd0;
  assign decode_speculative            = 1'd1;
  assign equals_units$000$clk          = clk;
  assign equals_units$000$compare_in_a = decode_inst[6:0];
  assign equals_units$000$compare_in_b = 7'd99;
  assign equals_units$000$reset        = reset;
  assign gen_data                      = lookup_out;
  assign gen_inst                      = decode_inst;
  assign lookup_out                    = lut$lookup_out;
  assign lut$clk                       = clk;
  assign lut$lookup_in_[2:0]           = decode_inst[14:12];
  assign lut$reset                     = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_result(rs=result_field_slice.start, re=result_field_slice.stop):
  //       s.decode_result.v = 0
  //       s.decode_result[rs:re].v = s.gen_payload

  // logic for connect_result()
  always @ (*) begin
    decode_result = 0;
    decode_result[(3)-1:0] = gen_payload;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_success():
  //       s.decode_success.v = s.gen_valid & s.and_unit.op_out

  // logic for compute_success()
  always @ (*) begin
    decode_success = (gen_valid&and_unit$op_out);
  end


endmodule // GenDecoder_0x687c848ae02befc7

//-----------------------------------------------------------------------------
// LookupTable_0x7098a106e042a7dc
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(3)) -> (valid: Bits(1), out: Bits(3))", "mapping": {"0": "type_=0x0:unsigned=0x0", "1": "type_=0x1:unsigned=0x0", "4": "type_=0x2:unsigned=0x0", "5": "type_=0x3:unsigned=0x0", "6": "type_=0x2:unsigned=0x1", "7": "type_=0x3:unsigned=0x1"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0x7098a106e042a7dc
(
  input  logic [   0:0] clk,
  input  logic [   2:0] lookup_in_,
  output logic [   2:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   2:0] mux$mux_default;
  logic   [   2:0] mux$mux_in_$000;
  logic   [   2:0] mux$mux_in_$001;
  logic   [   2:0] mux$mux_in_$002;
  logic   [   2:0] mux$mux_in_$003;
  logic   [   2:0] mux$mux_in_$004;
  logic   [   2:0] mux$mux_in_$005;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   2:0] mux$mux_select;
  logic   [   2:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x49a70fe32bf90ddf mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .mux_in_$003 ( mux$mux_in_$003 ),
    .mux_in_$004 ( mux$mux_in_$004 ),
    .mux_in_$005 ( mux$mux_in_$005 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 3'd0;
  assign mux$mux_in_$000 = 3'd0;
  assign mux$mux_in_$001 = 3'd1;
  assign mux$mux_in_$002 = 3'd2;
  assign mux$mux_in_$003 = 3'd3;
  assign mux$mux_in_$004 = 3'd6;
  assign mux$mux_in_$005 = 3'd7;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0x7098a106e042a7dc

//-----------------------------------------------------------------------------
// CaseMux_0x49a70fe32bf90ddf
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(3), in_: Bits(3) [6], select: Bits(3)) -> (out: Bits(3), matched: Bits(1))", "svalues": ["0", "1", "4", "5", "6", "7"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x49a70fe32bf90ddf
(
  input  logic [   0:0] clk,
  input  logic [   2:0] mux_default,
  input  logic [   2:0] mux_in_$000,
  input  logic [   2:0] mux_in_$001,
  input  logic [   2:0] mux_in_$002,
  input  logic [   2:0] mux_in_$003,
  input  logic [   2:0] mux_in_$004,
  input  logic [   2:0] mux_in_$005,
  output logic [   0:0] mux_matched,
  output logic [   2:0] mux_out,
  input  logic [   2:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   2:0] out_chain$000;
  logic   [   2:0] out_chain$001;
  logic   [   2:0] out_chain$002;
  logic   [   2:0] out_chain$003;
  logic   [   2:0] out_chain$004;
  logic   [   2:0] out_chain$005;
  logic   [   2:0] out_chain$006;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;
  logic   [   0:0] valid_chain$003;
  logic   [   0:0] valid_chain$004;
  logic   [   0:0] valid_chain$005;
  logic   [   0:0] valid_chain$006;


  // signal connections
  assign mux_matched     = valid_chain$006;
  assign mux_out         = out_chain$006;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   2:0] mux_in_[0:5];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  assign mux_in_[  3] = mux_in_$003;
  assign mux_in_[  4] = mux_in_$004;
  assign mux_in_[  5] = mux_in_$005;
  logic    [   2:0] out_chain[0:6];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  assign out_chain$003 = out_chain[  3];
  assign out_chain$004 = out_chain[  4];
  assign out_chain$005 = out_chain[  5];
  assign out_chain$006 = out_chain[  6];
  logic    [   0:0] valid_chain[0:6];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];
  assign valid_chain$003 = valid_chain[  3];
  assign valid_chain$004 = valid_chain[  4];
  assign valid_chain$005 = valid_chain[  5];
  assign valid_chain$006 = valid_chain[  6];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 0)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 1)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 4)) begin
      out_chain[3] = mux_in_[2];
      valid_chain[3] = 1;
    end
    else begin
      out_chain[3] = out_chain[2];
      valid_chain[3] = valid_chain[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 5)) begin
      out_chain[4] = mux_in_[3];
      valid_chain[4] = 1;
    end
    else begin
      out_chain[4] = out_chain[3];
      valid_chain[4] = valid_chain[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 6)) begin
      out_chain[5] = mux_in_[4];
      valid_chain[5] = 1;
    end
    else begin
      out_chain[5] = out_chain[4];
      valid_chain[5] = valid_chain[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 7)) begin
      out_chain[6] = mux_in_[5];
      valid_chain[6] = 1;
    end
    else begin
      out_chain[6] = out_chain[5];
      valid_chain[6] = valid_chain[5];
    end
  end


endmodule // CaseMux_0x49a70fe32bf90ddf

//-----------------------------------------------------------------------------
// ImmDecoder_0x67749655d31303e2
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.imm_decoder {"interface": "decode (type_: Bits(3), inst: Bits(32)) -> (imm: Bits(21))"}
// PyMTL: verilator_xinit = zeros
module ImmDecoder_0x67749655d31303e2
(
  input  logic [   0:0] clk,
  output logic [  20:0] decode_imm,
  input  logic [  31:0] decode_inst,
  input  logic [   2:0] decode_type_,
  input  logic [   0:0] reset
);

  // register declarations
  logic    [  12:0] imm_b;
  logic    [   4:0] imm_c;
  logic    [  11:0] imm_i;
  logic    [  20:0] imm_j;
  logic    [  11:0] imm_s;
  logic    [   4:0] imm_shamt32;
  logic    [   5:0] imm_shamt64;
  logic    [  19:0] imm_u;

  // localparam declarations
  localparam IMM_TYPE_B = 3'd2;
  localparam IMM_TYPE_C = 3'd5;
  localparam IMM_TYPE_I = 3'd0;
  localparam IMM_TYPE_J = 3'd4;
  localparam IMM_TYPE_S = 3'd1;
  localparam IMM_TYPE_SHAMT32 = 3'd6;
  localparam IMM_TYPE_SHAMT64 = 3'd7;
  localparam IMM_TYPE_U = 3'd3;
  localparam imm_len = 21;

  // mux temporaries
  logic   [  20:0] mux$mux_in_$000;
  logic   [  20:0] mux$mux_in_$001;
  logic   [  20:0] mux$mux_in_$002;
  logic   [  20:0] mux$mux_in_$003;
  logic   [  20:0] mux$mux_in_$004;
  logic   [  20:0] mux$mux_in_$005;
  logic   [  20:0] mux$mux_in_$006;
  logic   [  20:0] mux$mux_in_$007;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   2:0] mux$mux_select;
  logic   [  20:0] mux$mux_out;

  Mux_0x677626a735201326 mux
  (
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .mux_in_$003 ( mux$mux_in_$003 ),
    .mux_in_$004 ( mux$mux_in_$004 ),
    .mux_in_$005 ( mux$mux_in_$005 ),
    .mux_in_$006 ( mux$mux_in_$006 ),
    .mux_in_$007 ( mux$mux_in_$007 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out )
  );

  // signal connections
  assign decode_imm     = mux$mux_out;
  assign mux$clk        = clk;
  assign mux$mux_select = decode_type_;
  assign mux$reset      = reset;

  // array declarations
  logic    [  20:0] mux$mux_in_[0:7];
  assign mux$mux_in_$000 = mux$mux_in_[  0];
  assign mux$mux_in_$001 = mux$mux_in_[  1];
  assign mux$mux_in_$002 = mux$mux_in_[  2];
  assign mux$mux_in_$003 = mux$mux_in_[  3];
  assign mux$mux_in_$004 = mux$mux_in_[  4];
  assign mux$mux_in_$005 = mux$mux_in_[  5];
  assign mux$mux_in_$006 = mux$mux_in_[  6];
  assign mux$mux_in_$007 = mux$mux_in_[  7];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_imm():
  //       s.imm_i.v = s.decode_inst.i_imm
  //       s.imm_s.v = concat(s.decode_inst.s_imm1, s.decode_inst.s_imm0)
  //       s.imm_b.v = (
  //           concat(s.decode_inst.b_imm3, s.decode_inst.b_imm2,
  //                  s.decode_inst.b_imm1, s.decode_inst.b_imm0, Bits(1, 0)))
  //       s.imm_u.v = s.decode_inst.u_imm
  //       s.imm_j.v = concat(s.decode_inst.j_imm3, s.decode_inst.j_imm2,
  //                          s.decode_inst.j_imm1, s.decode_inst.j_imm0, Bits(1, 0))
  //       s.imm_c.v = s.decode_inst.c_imm
  //       s.imm_shamt32.v = s.decode_inst.shamt32
  //       s.imm_shamt64.v = s.decode_inst.shamt64
  //
  //       s.mux.mux_in_[ImmType.IMM_TYPE_I].v = sext(s.imm_i, imm_len)
  //       s.mux.mux_in_[ImmType.IMM_TYPE_S].v = sext(s.imm_s, imm_len)
  //       s.mux.mux_in_[ImmType.IMM_TYPE_B].v = sext(s.imm_b, imm_len)
  //       s.mux.mux_in_[ImmType.IMM_TYPE_U].v = sext(s.imm_u, imm_len)
  //       s.mux.mux_in_[ImmType.IMM_TYPE_J].v = sext(s.imm_j, imm_len)
  //       s.mux.mux_in_[ImmType.IMM_TYPE_C].v = zext(s.imm_c, imm_len)
  //       s.mux.mux_in_[ImmType.IMM_TYPE_SHAMT32].v = zext(s.imm_shamt32, imm_len)
  //       s.mux.mux_in_[ImmType.IMM_TYPE_SHAMT64].v = zext(s.imm_shamt64, imm_len)

  // logic for handle_imm()
  always @ (*) begin
    imm_i = decode_inst[(32)-1:20];
    imm_s = { decode_inst[(32)-1:25],decode_inst[(12)-1:7] };
    imm_b = { decode_inst[(32)-1:31],decode_inst[(8)-1:7],decode_inst[(31)-1:25],decode_inst[(12)-1:8],1'd0 };
    imm_u = decode_inst[(32)-1:12];
    imm_j = { decode_inst[(32)-1:31],decode_inst[(20)-1:12],decode_inst[(21)-1:20],decode_inst[(31)-1:21],1'd0 };
    imm_c = decode_inst[(20)-1:15];
    imm_shamt32 = decode_inst[(25)-1:20];
    imm_shamt64 = decode_inst[(26)-1:20];
    mux$mux_in_[IMM_TYPE_I] = { { imm_len-12 { imm_i[11] } }, imm_i };
    mux$mux_in_[IMM_TYPE_S] = { { imm_len-12 { imm_s[11] } }, imm_s };
    mux$mux_in_[IMM_TYPE_B] = { { imm_len-13 { imm_b[12] } }, imm_b };
    mux$mux_in_[IMM_TYPE_U] = { { imm_len-20 { imm_u[19] } }, imm_u };
    mux$mux_in_[IMM_TYPE_J] = { { imm_len-21 { imm_j[20] } }, imm_j };
    mux$mux_in_[IMM_TYPE_C] = { { imm_len-5 { 1'b0 } }, imm_c };
    mux$mux_in_[IMM_TYPE_SHAMT32] = { { imm_len-5 { 1'b0 } }, imm_shamt32 };
    mux$mux_in_[IMM_TYPE_SHAMT64] = { { imm_len-6 { 1'b0 } }, imm_shamt64 };
  end


endmodule // ImmDecoder_0x67749655d31303e2

//-----------------------------------------------------------------------------
// Mux_0x677626a735201326
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.mux {"dtype": 21, "nports": 8}
// PyMTL: verilator_xinit = zeros
module Mux_0x677626a735201326
(
  input  logic [   0:0] clk,
  input  logic [  20:0] mux_in_$000,
  input  logic [  20:0] mux_in_$001,
  input  logic [  20:0] mux_in_$002,
  input  logic [  20:0] mux_in_$003,
  input  logic [  20:0] mux_in_$004,
  input  logic [  20:0] mux_in_$005,
  input  logic [  20:0] mux_in_$006,
  input  logic [  20:0] mux_in_$007,
  output logic  [  20:0] mux_out,
  input  logic [   2:0] mux_select,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nports = 8;


  // array declarations
  logic   [  20:0] mux_in_[0:7];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  assign mux_in_[  3] = mux_in_$003;
  assign mux_in_[  4] = mux_in_$004;
  assign mux_in_[  5] = mux_in_$005;
  assign mux_in_[  6] = mux_in_$006;
  assign mux_in_[  7] = mux_in_$007;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def select():
  //       assert s.mux_select < nports
  //       s.mux_out.v = s.mux_in_[s.mux_select]

  // logic for select()
  always @ (*) begin
    mux_out = mux_in_[mux_select];
  end


endmodule // Mux_0x677626a735201326

//-----------------------------------------------------------------------------
// GS11LBranchStage20LBranchDropController_0xc628584b4321be9
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"args": ["process <C> (in_: Bits(251)) -> (accepted: Bits(1), out: Bits(146))"], "kwargs": {}}
// PyMTL: verilator_xinit = zeros
module GS11LBranchStage20LBranchDropController_0xc628584b4321be9
(
  output logic [   0:0] cflow_redirect_call,
  output logic [   0:0] cflow_redirect_force,
  output logic [   3:0] cflow_redirect_seq,
  output logic [   0:0] cflow_redirect_spec_idx,
  output logic [  63:0] cflow_redirect_target,
  input  logic [   0:0] clk,
  input  logic [ 250:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 145:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // pipeline_stage temporaries
  logic   [   0:0] pipeline_stage$check_keep;
  logic   [ 250:0] pipeline_stage$in_peek_msg;
  logic   [   0:0] pipeline_stage$clk;
  logic   [   4:0] pipeline_stage$kill_notify_msg;
  logic   [   0:0] pipeline_stage$in_peek_rdy;
  logic   [   0:0] pipeline_stage$process_accepted;
  logic   [ 145:0] pipeline_stage$check_out;
  logic   [   0:0] pipeline_stage$reset;
  logic   [ 145:0] pipeline_stage$process_out;
  logic   [   0:0] pipeline_stage$take_call;
  logic   [   0:0] pipeline_stage$process_call;
  logic   [ 145:0] pipeline_stage$check_in_;
  logic   [ 145:0] pipeline_stage$peek_msg;
  logic   [   4:0] pipeline_stage$check_msg;
  logic   [   0:0] pipeline_stage$in_take_call;
  logic   [   0:0] pipeline_stage$peek_rdy;
  logic   [ 250:0] pipeline_stage$process_in_;

  PipelineStage_0x3bdbe2fe9599a701 pipeline_stage
  (
    .check_keep       ( pipeline_stage$check_keep ),
    .in_peek_msg      ( pipeline_stage$in_peek_msg ),
    .clk              ( pipeline_stage$clk ),
    .kill_notify_msg  ( pipeline_stage$kill_notify_msg ),
    .in_peek_rdy      ( pipeline_stage$in_peek_rdy ),
    .process_accepted ( pipeline_stage$process_accepted ),
    .check_out        ( pipeline_stage$check_out ),
    .reset            ( pipeline_stage$reset ),
    .process_out      ( pipeline_stage$process_out ),
    .take_call        ( pipeline_stage$take_call ),
    .process_call     ( pipeline_stage$process_call ),
    .check_in_        ( pipeline_stage$check_in_ ),
    .peek_msg         ( pipeline_stage$peek_msg ),
    .check_msg        ( pipeline_stage$check_msg ),
    .in_take_call     ( pipeline_stage$in_take_call ),
    .peek_rdy         ( pipeline_stage$peek_rdy ),
    .process_in_      ( pipeline_stage$process_in_ )
  );

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [ 145:0] drop_controller$check_in_;
  logic   [   4:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [ 145:0] drop_controller$check_out;

  PipelineKillDropController_0x52612c5d4a64ec3 drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // stage temporaries
  logic   [   0:0] stage$process_call;
  logic   [   0:0] stage$clk;
  logic   [   0:0] stage$reset;
  logic   [ 250:0] stage$process_in_;
  logic   [   0:0] stage$cflow_redirect_call;
  logic   [   0:0] stage$process_accepted;
  logic   [  63:0] stage$cflow_redirect_target;
  logic   [   3:0] stage$cflow_redirect_seq;
  logic   [   0:0] stage$cflow_redirect_force;
  logic   [ 145:0] stage$process_out;
  logic   [   0:0] stage$cflow_redirect_spec_idx;

  BranchStage_0x5126114ec6ac2c47 stage
  (
    .process_call            ( stage$process_call ),
    .clk                     ( stage$clk ),
    .reset                   ( stage$reset ),
    .process_in_             ( stage$process_in_ ),
    .cflow_redirect_call     ( stage$cflow_redirect_call ),
    .process_accepted        ( stage$process_accepted ),
    .cflow_redirect_target   ( stage$cflow_redirect_target ),
    .cflow_redirect_seq      ( stage$cflow_redirect_seq ),
    .cflow_redirect_force    ( stage$cflow_redirect_force ),
    .process_out             ( stage$process_out ),
    .cflow_redirect_spec_idx ( stage$cflow_redirect_spec_idx )
  );

  // signal connections
  assign cflow_redirect_call             = stage$cflow_redirect_call;
  assign cflow_redirect_force            = stage$cflow_redirect_force;
  assign cflow_redirect_seq              = stage$cflow_redirect_seq;
  assign cflow_redirect_spec_idx         = stage$cflow_redirect_spec_idx;
  assign cflow_redirect_target           = stage$cflow_redirect_target;
  assign drop_controller$check_in_       = pipeline_stage$check_in_;
  assign drop_controller$check_msg       = pipeline_stage$check_msg;
  assign drop_controller$clk             = clk;
  assign drop_controller$reset           = reset;
  assign in_take_call                    = pipeline_stage$in_take_call;
  assign peek_msg                        = pipeline_stage$peek_msg;
  assign peek_rdy                        = pipeline_stage$peek_rdy;
  assign pipeline_stage$check_keep       = drop_controller$check_keep;
  assign pipeline_stage$check_out        = drop_controller$check_out;
  assign pipeline_stage$clk              = clk;
  assign pipeline_stage$in_peek_msg      = in_peek_msg;
  assign pipeline_stage$in_peek_rdy      = in_peek_rdy;
  assign pipeline_stage$kill_notify_msg  = kill_notify_msg;
  assign pipeline_stage$process_accepted = stage$process_accepted;
  assign pipeline_stage$process_out      = stage$process_out;
  assign pipeline_stage$reset            = reset;
  assign pipeline_stage$take_call        = take_call;
  assign stage$clk                       = clk;
  assign stage$process_call              = pipeline_stage$process_call;
  assign stage$process_in_               = pipeline_stage$process_in_;
  assign stage$reset                     = reset;



endmodule // GS11LBranchStage20LBranchDropController_0xc628584b4321be9

//-----------------------------------------------------------------------------
// BranchStage_0x5126114ec6ac2c47
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.backend.branch {"branch_interface": "process <C> (in_: Bits(251)) -> (accepted: Bits(1), out: Bits(146))"}
// PyMTL: verilator_xinit = zeros
module BranchStage_0x5126114ec6ac2c47
(
  output logic [   0:0] cflow_redirect_call,
  output logic [   0:0] cflow_redirect_force,
  output logic [   3:0] cflow_redirect_seq,
  output logic [   0:0] cflow_redirect_spec_idx,
  output logic [  63:0] cflow_redirect_target,
  input  logic [   0:0] clk,
  output logic [   0:0] process_accepted,
  input  logic [   0:0] process_call,
  input  logic [ 250:0] process_in_,
  output logic  [ 145:0] process_out,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [ 250:0] msg_;


  // register declarations
  logic    [  63:0] branch_target_;
  logic    [  63:0] imm_;
  logic    [  20:0] msg_imm_;
  logic    [   0:0] take_branch_;

  // localparam declarations
  localparam data_len = 64;

  // op_lut_ temporaries
  logic   [   0:0] op_lut_$clk;
  logic   [   0:0] op_lut_$reset;
  logic   [   1:0] op_lut_$lookup_in_;
  logic   [   1:0] op_lut_$lookup_out;
  logic   [   0:0] op_lut_$lookup_valid;

  LookupTable_0x4b32e275e4f79d2a op_lut_
  (
    .clk          ( op_lut_$clk ),
    .reset        ( op_lut_$reset ),
    .lookup_in_   ( op_lut_$lookup_in_ ),
    .lookup_out   ( op_lut_$lookup_out ),
    .lookup_valid ( op_lut_$lookup_valid )
  );

  // cmp_ temporaries
  logic   [   0:0] cmp_$exec_unsigned;
  logic   [   0:0] cmp_$clk;
  logic   [  63:0] cmp_$exec_src1;
  logic   [  63:0] cmp_$exec_src0;
  logic   [   1:0] cmp_$exec_func;
  logic   [   0:0] cmp_$exec_call;
  logic   [   0:0] cmp_$reset;
  logic   [   0:0] cmp_$exec_res;
  logic   [   0:0] cmp_$exec_rdy;

  Comparator_0x53ba82e9f98ca135 cmp_
  (
    .exec_unsigned ( cmp_$exec_unsigned ),
    .clk           ( cmp_$clk ),
    .exec_src1     ( cmp_$exec_src1 ),
    .exec_src0     ( cmp_$exec_src0 ),
    .exec_func     ( cmp_$exec_func ),
    .exec_call     ( cmp_$exec_call ),
    .reset         ( cmp_$reset ),
    .exec_res      ( cmp_$exec_res ),
    .exec_rdy      ( cmp_$exec_rdy )
  );

  // signal connections
  assign cflow_redirect_call     = process_call;
  assign cflow_redirect_force    = 1'd0;
  assign cflow_redirect_seq      = msg_[69:66];
  assign cflow_redirect_spec_idx = msg_[71:71];
  assign cflow_redirect_target   = branch_target_;
  assign cmp_$clk                = clk;
  assign cmp_$exec_call          = process_call;
  assign cmp_$exec_func          = op_lut_$lookup_out;
  assign cmp_$exec_src0          = msg_[138:75];
  assign cmp_$exec_src1          = msg_[203:140];
  assign cmp_$exec_unsigned      = msg_[238:238];
  assign cmp_$reset              = reset;
  assign msg_                    = process_in_;
  assign op_lut_$clk             = clk;
  assign op_lut_$lookup_in_      = msg_[237:236];
  assign op_lut_$reset           = reset;
  assign process_accepted        = 1'd1;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_take_branch():
  //       s.take_branch_.v = 0
  //       # TODO handle branches that are not conditional
  //       s.take_branch_.v = s.cmp_.exec_res

  // logic for set_take_branch()
  always @ (*) begin
    take_branch_ = 0;
    take_branch_ = cmp_$exec_res;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_target():
  //       s.msg_imm_.v = s.msg_.imm
  //       # PYMTL_BROKEN: sext(s.msg_.imm) does not create valid verilog
  //       # Vivado errors: "range is not allowed in prefix"
  //       s.imm_.v = sext(s.msg_imm_, data_len)
  //       if s.take_branch_:
  //         s.branch_target_.v = s.msg_.hdr_pc + s.imm_
  //       else:
  //         s.branch_target_.v = s.msg_.hdr_pc + 4

  // logic for compute_target()
  always @ (*) begin
    msg_imm_ = msg_[(233)-1:212];
    imm_ = { { data_len-21 { msg_imm_[20] } }, msg_imm_ };
    if (take_branch_) begin
      branch_target_ = (msg_[(66)-1:2]+imm_);
    end
    else begin
      branch_target_ = (msg_[(66)-1:2]+4);
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_value_reg_input():
  //       s.process_out.v = 0
  //       s.process_out.hdr.v = s.msg_.hdr

  // logic for set_value_reg_input()
  always @ (*) begin
    process_out = 0;
    process_out[(74)-1:0] = msg_[(74)-1:0];
  end


endmodule // BranchStage_0x5126114ec6ac2c47

//-----------------------------------------------------------------------------
// LookupTable_0x4b32e275e4f79d2a
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.lookup_table {"interface": "lookup (in_: Bits(2)) -> (valid: Bits(1), out: Bits(2))", "mapping": {"0": "0", "1": "1", "2": "2", "3": "3"}}
// PyMTL: verilator_xinit = zeros
module LookupTable_0x4b32e275e4f79d2a
(
  input  logic [   0:0] clk,
  input  logic [   1:0] lookup_in_,
  output logic [   1:0] lookup_out,
  output logic [   0:0] lookup_valid,
  input  logic [   0:0] reset
);

  // mux temporaries
  logic   [   1:0] mux$mux_default;
  logic   [   1:0] mux$mux_in_$000;
  logic   [   1:0] mux$mux_in_$001;
  logic   [   1:0] mux$mux_in_$002;
  logic   [   1:0] mux$mux_in_$003;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   1:0] mux$mux_select;
  logic   [   1:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x4d0f7376ef889108 mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .mux_in_$003 ( mux$mux_in_$003 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign lookup_out      = mux$mux_out;
  assign lookup_valid    = mux$mux_matched;
  assign mux$clk         = clk;
  assign mux$mux_default = 2'd0;
  assign mux$mux_in_$000 = 2'd0;
  assign mux$mux_in_$001 = 2'd1;
  assign mux$mux_in_$002 = 2'd2;
  assign mux$mux_in_$003 = 2'd3;
  assign mux$mux_select  = lookup_in_;
  assign mux$reset       = reset;



endmodule // LookupTable_0x4b32e275e4f79d2a

//-----------------------------------------------------------------------------
// CaseMux_0x4d0f7376ef889108
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(2), in_: Bits(2) [4], select: Bits(2)) -> (out: Bits(2), matched: Bits(1))", "svalues": ["0", "1", "2", "3"]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x4d0f7376ef889108
(
  input  logic [   0:0] clk,
  input  logic [   1:0] mux_default,
  input  logic [   1:0] mux_in_$000,
  input  logic [   1:0] mux_in_$001,
  input  logic [   1:0] mux_in_$002,
  input  logic [   1:0] mux_in_$003,
  output logic [   0:0] mux_matched,
  output logic [   1:0] mux_out,
  input  logic [   1:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   1:0] out_chain$000;
  logic   [   1:0] out_chain$001;
  logic   [   1:0] out_chain$002;
  logic   [   1:0] out_chain$003;
  logic   [   1:0] out_chain$004;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;
  logic   [   0:0] valid_chain$003;
  logic   [   0:0] valid_chain$004;


  // signal connections
  assign mux_matched     = valid_chain$004;
  assign mux_out         = out_chain$004;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [   1:0] mux_in_[0:3];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  assign mux_in_[  3] = mux_in_$003;
  logic    [   1:0] out_chain[0:4];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  assign out_chain$003 = out_chain[  3];
  assign out_chain$004 = out_chain[  4];
  logic    [   0:0] valid_chain[0:4];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];
  assign valid_chain$003 = valid_chain[  3];
  assign valid_chain$004 = valid_chain[  4];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 0)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 1)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 2)) begin
      out_chain[3] = mux_in_[2];
      valid_chain[3] = 1;
    end
    else begin
      out_chain[3] = out_chain[2];
      valid_chain[3] = valid_chain[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 3)) begin
      out_chain[4] = mux_in_[3];
      valid_chain[4] = 1;
    end
    else begin
      out_chain[4] = out_chain[3];
      valid_chain[4] = valid_chain[3];
    end
  end


endmodule // CaseMux_0x4d0f7376ef889108

//-----------------------------------------------------------------------------
// Comparator_0x53ba82e9f98ca135
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.comparator {"alu_interface": "exec <CR> (src0: Bits(64), src1: Bits(64), unsigned: Bits(1), func: Bits(2)) -> (res: Bits(1))"}
// PyMTL: verilator_xinit = zeros
module Comparator_0x53ba82e9f98ca135
(
  input  logic [   0:0] clk,
  input  logic [   0:0] exec_call,
  input  logic [   1:0] exec_func,
  output logic [   0:0] exec_rdy,
  output logic [   0:0] exec_res,
  input  logic [  63:0] exec_src0,
  input  logic [  63:0] exec_src1,
  input  logic [   0:0] exec_unsigned,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   1:0] func_;


  // register declarations
  logic    [   0:0] eq_;
  logic    [   0:0] lt_;
  logic    [   0:0] res_;
  logic    [  63:0] s0_;
  logic    [  62:0] s0_lower_;
  logic    [   0:0] s0_up_;
  logic    [  63:0] s1_;
  logic    [  62:0] s1_lower_;
  logic    [   0:0] s1_up_;

  // localparam declarations
  localparam CMP_EQ = 2'd0;
  localparam CMP_GE = 2'd3;
  localparam CMP_LT = 2'd2;
  localparam CMP_NE = 2'd1;
  localparam XLEN_M1 = 63;

  // signal connections
  assign exec_rdy = 1'd1;
  assign exec_res = res_;
  assign func_    = exec_func;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_flags():
  //       s.eq_.v = s.s0_ == s.s1_
  //       s.lt_.v = s.s0_ < s.s1_

  // logic for set_flags()
  always @ (*) begin
    eq_ = (s0_ == s1_);
    lt_ = (s0_ < s1_);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_signed():
  //       # We flip the upper most bit if signed
  //       s.s0_up_.v = s.exec_src0[
  //           XLEN_M1] if s.exec_unsigned else not s.exec_src0[XLEN_M1]
  //       s.s1_up_.v = s.exec_src1[
  //           XLEN_M1] if s.exec_unsigned else not s.exec_src1[XLEN_M1]
  //       s.s0_lower_.v = s.exec_src0[0:XLEN_M1]
  //       s.s1_lower_.v = s.exec_src1[0:XLEN_M1]
  //       # Now we can concat and compare
  //       s.s0_.v = concat(s.s0_up_, s.s0_lower_)
  //       s.s1_.v = concat(s.s1_up_, s.s1_lower_)

  // logic for set_signed()
  always @ (*) begin
    s0_up_ = exec_unsigned ? exec_src0[XLEN_M1] : !exec_src0[XLEN_M1];
    s1_up_ = exec_unsigned ? exec_src1[XLEN_M1] : !exec_src1[XLEN_M1];
    s0_lower_ = exec_src0[(XLEN_M1)-1:0];
    s1_lower_ = exec_src1[(XLEN_M1)-1:0];
    s0_ = { s0_up_,s0_lower_ };
    s1_ = { s1_up_,s1_lower_ };
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def eval_comb():
  //       s.res_.v = 0
  //       if s.exec_call:
  //         if s.func_ == CMPFunc.CMP_EQ:
  //           s.res_.v = s.eq_
  //         elif s.func_ == CMPFunc.CMP_NE:
  //           s.res_.v = not s.eq_
  //         elif s.func_ == CMPFunc.CMP_LT:
  //           s.res_.v = s.lt_
  //         elif s.func_ == CMPFunc.CMP_GE:
  //           s.res_.v = not s.lt_ or s.eq_

  // logic for eval_comb()
  always @ (*) begin
    res_ = 0;
    if (exec_call) begin
      if ((func_ == CMP_EQ)) begin
        res_ = eq_;
      end
      else begin
        if ((func_ == CMP_NE)) begin
          res_ = !eq_;
        end
        else begin
          if ((func_ == CMP_LT)) begin
            res_ = lt_;
          end
          else begin
            if ((func_ == CMP_GE)) begin
              res_ = (!lt_||eq_);
            end
            else begin
            end
          end
        end
      end
    end
    else begin
    end
  end


endmodule // Comparator_0x53ba82e9f98ca135

//-----------------------------------------------------------------------------
// GS8LCSRStage17LCSRDropController_0xc628584b4321be9
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"args": ["process <C> (in_: Bits(251)) -> (accepted: Bits(1), out: Bits(146))"], "kwargs": {}}
// PyMTL: verilator_xinit = zeros
module GS8LCSRStage17LCSRDropController_0xc628584b4321be9
(
  input  logic [   0:0] clk,
  output logic [   0:0] csr_op_call,
  output logic [  11:0] csr_op_csr,
  input  logic [  63:0] csr_op_old,
  output logic [   1:0] csr_op_op,
  output logic [   0:0] csr_op_rs1_is_x0,
  input  logic [   0:0] csr_op_success,
  output logic [  63:0] csr_op_value,
  input  logic [ 250:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 145:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // pipeline_stage temporaries
  logic   [   0:0] pipeline_stage$check_keep;
  logic   [ 250:0] pipeline_stage$in_peek_msg;
  logic   [   0:0] pipeline_stage$clk;
  logic   [   4:0] pipeline_stage$kill_notify_msg;
  logic   [   0:0] pipeline_stage$in_peek_rdy;
  logic   [   0:0] pipeline_stage$process_accepted;
  logic   [ 145:0] pipeline_stage$check_out;
  logic   [   0:0] pipeline_stage$reset;
  logic   [ 145:0] pipeline_stage$process_out;
  logic   [   0:0] pipeline_stage$take_call;
  logic   [   0:0] pipeline_stage$process_call;
  logic   [ 145:0] pipeline_stage$check_in_;
  logic   [ 145:0] pipeline_stage$peek_msg;
  logic   [   4:0] pipeline_stage$check_msg;
  logic   [   0:0] pipeline_stage$in_take_call;
  logic   [   0:0] pipeline_stage$peek_rdy;
  logic   [ 250:0] pipeline_stage$process_in_;

  PipelineStage_0x3bdbe2fe9599a701 pipeline_stage
  (
    .check_keep       ( pipeline_stage$check_keep ),
    .in_peek_msg      ( pipeline_stage$in_peek_msg ),
    .clk              ( pipeline_stage$clk ),
    .kill_notify_msg  ( pipeline_stage$kill_notify_msg ),
    .in_peek_rdy      ( pipeline_stage$in_peek_rdy ),
    .process_accepted ( pipeline_stage$process_accepted ),
    .check_out        ( pipeline_stage$check_out ),
    .reset            ( pipeline_stage$reset ),
    .process_out      ( pipeline_stage$process_out ),
    .take_call        ( pipeline_stage$take_call ),
    .process_call     ( pipeline_stage$process_call ),
    .check_in_        ( pipeline_stage$check_in_ ),
    .peek_msg         ( pipeline_stage$peek_msg ),
    .check_msg        ( pipeline_stage$check_msg ),
    .in_take_call     ( pipeline_stage$in_take_call ),
    .peek_rdy         ( pipeline_stage$peek_rdy ),
    .process_in_      ( pipeline_stage$process_in_ )
  );

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [ 145:0] drop_controller$check_in_;
  logic   [   4:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [ 145:0] drop_controller$check_out;

  PipelineKillDropController_0x52612c5d4a64ec3 drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // stage temporaries
  logic   [   0:0] stage$process_call;
  logic   [   0:0] stage$csr_op_success;
  logic   [  63:0] stage$csr_op_old;
  logic   [   0:0] stage$clk;
  logic   [   0:0] stage$reset;
  logic   [ 250:0] stage$process_in_;
  logic   [   1:0] stage$csr_op_op;
  logic   [   0:0] stage$csr_op_call;
  logic   [   0:0] stage$process_accepted;
  logic   [   0:0] stage$csr_op_rs1_is_x0;
  logic   [  11:0] stage$csr_op_csr;
  logic   [  63:0] stage$csr_op_value;
  logic   [ 145:0] stage$process_out;

  CSRStage_0x2aafa7618480546 stage
  (
    .process_call     ( stage$process_call ),
    .csr_op_success   ( stage$csr_op_success ),
    .csr_op_old       ( stage$csr_op_old ),
    .clk              ( stage$clk ),
    .reset            ( stage$reset ),
    .process_in_      ( stage$process_in_ ),
    .csr_op_op        ( stage$csr_op_op ),
    .csr_op_call      ( stage$csr_op_call ),
    .process_accepted ( stage$process_accepted ),
    .csr_op_rs1_is_x0 ( stage$csr_op_rs1_is_x0 ),
    .csr_op_csr       ( stage$csr_op_csr ),
    .csr_op_value     ( stage$csr_op_value ),
    .process_out      ( stage$process_out )
  );

  // signal connections
  assign csr_op_call                     = stage$csr_op_call;
  assign csr_op_csr                      = stage$csr_op_csr;
  assign csr_op_op                       = stage$csr_op_op;
  assign csr_op_rs1_is_x0                = stage$csr_op_rs1_is_x0;
  assign csr_op_value                    = stage$csr_op_value;
  assign drop_controller$check_in_       = pipeline_stage$check_in_;
  assign drop_controller$check_msg       = pipeline_stage$check_msg;
  assign drop_controller$clk             = clk;
  assign drop_controller$reset           = reset;
  assign in_take_call                    = pipeline_stage$in_take_call;
  assign peek_msg                        = pipeline_stage$peek_msg;
  assign peek_rdy                        = pipeline_stage$peek_rdy;
  assign pipeline_stage$check_keep       = drop_controller$check_keep;
  assign pipeline_stage$check_out        = drop_controller$check_out;
  assign pipeline_stage$clk              = clk;
  assign pipeline_stage$in_peek_msg      = in_peek_msg;
  assign pipeline_stage$in_peek_rdy      = in_peek_rdy;
  assign pipeline_stage$kill_notify_msg  = kill_notify_msg;
  assign pipeline_stage$process_accepted = stage$process_accepted;
  assign pipeline_stage$process_out      = stage$process_out;
  assign pipeline_stage$reset            = reset;
  assign pipeline_stage$take_call        = take_call;
  assign stage$clk                       = clk;
  assign stage$csr_op_old                = csr_op_old;
  assign stage$csr_op_success            = csr_op_success;
  assign stage$process_call              = pipeline_stage$process_call;
  assign stage$process_in_               = pipeline_stage$process_in_;
  assign stage$reset                     = reset;



endmodule // GS8LCSRStage17LCSRDropController_0xc628584b4321be9

//-----------------------------------------------------------------------------
// CSRStage_0x2aafa7618480546
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.backend.csr {"interface": "process <C> (in_: Bits(251)) -> (accepted: Bits(1), out: Bits(146))"}
// PyMTL: verilator_xinit = zeros
module CSRStage_0x2aafa7618480546
(
  input  logic [   0:0] clk,
  output logic  [   0:0] csr_op_call,
  output logic  [  11:0] csr_op_csr,
  input  logic [  63:0] csr_op_old,
  output logic  [   1:0] csr_op_op,
  output logic  [   0:0] csr_op_rs1_is_x0,
  input  logic [   0:0] csr_op_success,
  output logic  [  63:0] csr_op_value,
  output logic [   0:0] process_accepted,
  input  logic [   0:0] process_call,
  input  logic [ 250:0] process_in_,
  output logic  [ 145:0] process_out,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam PIPELINE_MSG_STATUS_VALID = 2'd0;

  // signal connections
  assign process_accepted = 1'd1;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_process():
  //       s.process_out.v = 0
  //       s.process_out.hdr.v = s.process_in_.hdr
  //
  //       s.csr_op_csr.v = 0
  //       s.csr_op_op.v = 0
  //       s.csr_op_rs1_is_x0.v = 0
  //       s.csr_op_value.v = 0
  //       s.csr_op_call.v = 0
  //
  //       if s.process_call:
  //         if s.process_in_.hdr_status == PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID:
  //           s.process_out.rd_val_pair.v = s.process_in_.rd_val_pair
  //           s.process_out.result.v = s.csr_op_old
  //           s.csr_op_csr.v = s.process_in_.csr_msg_csr_num
  //           s.csr_op_op.v = s.process_in_.csr_msg_func
  //           s.csr_op_rs1_is_x0.v = s.process_in_.csr_msg_rs1_is_x0
  //           s.csr_op_value.v = s.process_in_.rs1
  //           s.csr_op_call.v = 1
  //
  //           # TODO handle failure
  //         else:
  //           s.process_out.exception_info.v = s.process_in_.exception_info

  // logic for handle_process()
  always @ (*) begin
    process_out = 0;
    process_out[(74)-1:0] = process_in_[(74)-1:0];
    csr_op_csr = 0;
    csr_op_op = 0;
    csr_op_rs1_is_x0 = 0;
    csr_op_value = 0;
    csr_op_call = 0;
    if (process_call) begin
      if ((process_in_[(2)-1:0] == PIPELINE_MSG_STATUS_VALID)) begin
        process_out[(81)-1:74] = process_in_[(211)-1:204];
        process_out[(146)-1:82] = csr_op_old;
        csr_op_csr = process_in_[(250)-1:238];
        csr_op_op = process_in_[(238)-1:236];
        csr_op_rs1_is_x0 = process_in_[(251)-1:250];
        csr_op_value = process_in_[(139)-1:75];
        csr_op_call = 1;
      end
      else begin
        process_out[(142)-1:74] = process_in_[(142)-1:74];
      end
    end
    else begin
    end
  end


endmodule // CSRStage_0x2aafa7618480546

//-----------------------------------------------------------------------------
// RedirectNotifier_0x76bce5ec03c6a79c
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.kill_unit {"xlen": 64}
// PyMTL: verilator_xinit = zeros
module RedirectNotifier_0x76bce5ec03c6a79c
(
  input  logic [   0:0] check_redirect_redirect,
  input  logic [  63:0] check_redirect_target,
  input  logic [   0:0] clk,
  output logic [   0:0] kill_notify_msg,
  input  logic [   0:0] reset
);

  // signal connections
  assign kill_notify_msg = check_redirect_redirect;



endmodule // RedirectNotifier_0x76bce5ec03c6a79c

//-----------------------------------------------------------------------------
// Issue_0x52678fcc1604a432
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.backend.issue {"interface": "kill_notify (msg: Bits(5)) -> (); peek <R> () -> (msg: Bits(142)); take <C> () -> ()", "num_pregs": 64, "num_slots": 2}
// PyMTL: verilator_xinit = zeros
module Issue_0x52678fcc1604a432
(
  input  logic [   0:0] clk,
  input  logic [  63:0] get_updated_mask,
  input  logic [ 141:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   0:0] is_ready_ready$000,
  input  logic [   0:0] is_ready_ready$001,
  output logic [   5:0] is_ready_tag$000,
  output logic [   5:0] is_ready_tag$001,
  input  logic [   4:0] kill_notify_msg,
  output logic  [ 141:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // logic declarations
  logic   [ 141:0] renamed_;


  // register declarations
  logic    [   0:0] accepted_;
  logic    [ 159:0] iq$add_value;
  logic    [ 141:0] iq_msg_in;
  logic    [ 159:0] iq_slot_in;

  // localparam declarations
  localparam PIPELINE_MSG_STATUS_VALID = 2'd0;

  // iq temporaries
  logic   [   0:0] iq$clk;
  logic   [   4:0] iq$kill_notify_msg;
  logic   [   5:0] iq$notify_value;
  logic   [   0:0] iq$reset;
  logic   [   0:0] iq$remove_call;
  logic   [   0:0] iq$notify_call;
  logic   [   0:0] iq$add_call;
  logic   [   0:0] iq$remove_rdy;
  logic   [   0:0] iq$add_rdy;
  logic   [ 159:0] iq$remove_value;

  CompactingIssueQueue_0x3a43583a53afd5b2 iq
  (
    .clk             ( iq$clk ),
    .kill_notify_msg ( iq$kill_notify_msg ),
    .notify_value    ( iq$notify_value ),
    .add_value       ( iq$add_value ),
    .reset           ( iq$reset ),
    .remove_call     ( iq$remove_call ),
    .notify_call     ( iq$notify_call ),
    .add_call        ( iq$add_call ),
    .remove_rdy      ( iq$remove_rdy ),
    .add_rdy         ( iq$add_rdy ),
    .remove_value    ( iq$remove_value )
  );

  // updated_ temporaries
  logic   [   0:0] updated_$clk;
  logic   [   0:0] updated_$reset;
  logic   [  63:0] updated_$decode_signal;
  logic   [   0:0] updated_$decode_valid;
  logic   [   5:0] updated_$decode_decoded;

  PriorityDecoder_0x2e5c0266b409153a updated_
  (
    .clk            ( updated_$clk ),
    .reset          ( updated_$reset ),
    .decode_signal  ( updated_$decode_signal ),
    .decode_valid   ( updated_$decode_valid ),
    .decode_decoded ( updated_$decode_decoded )
  );

  // signal connections
  assign in_take_call           = accepted_;
  assign iq$add_call            = accepted_;
  assign iq$clk                 = clk;
  assign iq$kill_notify_msg     = kill_notify_msg;
  assign iq$notify_call         = updated_$decode_valid;
  assign iq$notify_value        = updated_$decode_decoded;
  assign iq$remove_call         = take_call;
  assign iq$reset               = reset;
  assign is_ready_tag$000       = renamed_[80:75];
  assign is_ready_tag$001       = renamed_[87:82];
  assign peek_rdy               = iq$remove_rdy;
  assign renamed_               = in_peek_msg;
  assign updated_$clk           = clk;
  assign updated_$decode_signal = get_updated_mask;
  assign updated_$reset         = reset;

  // array declarations
  logic   [   0:0] is_ready_ready[0:1];
  assign is_ready_ready[  0] = is_ready_ready$000;
  assign is_ready_ready[  1] = is_ready_ready$001;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_accepted():
  //       s.accepted_.v = s.in_peek_rdy and s.iq.add_rdy

  // logic for set_accepted()
  always @ (*) begin
    accepted_ = (in_peek_rdy&&iq$add_rdy);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_input():
  //       s.iq_slot_in.v = 0
  //       # Copy header
  //       s.iq_msg_in.v = 0
  //       s.iq_msg_in.hdr.v = s.renamed_.hdr
  //       # Set the kill_opaque
  //       s.iq_slot_in.kill_opaque.v = s.renamed_.hdr_branch_mask
  //       # If there is an exception, make sure sources are invalid
  //       if s.renamed_.hdr_status != PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID:
  //         s.iq_slot_in.src0_val.v = 0
  //         s.iq_slot_in.src1_val.v = 0
  //         s.iq_msg_in.exception_info.v = s.renamed_.exception_info
  //       else:
  //         # Copy over the message contents
  //         s.iq_msg_in.execution_data.v = s.renamed_.execution_data
  //         s.iq_msg_in.rd.v = s.renamed_.rd
  //         s.iq_msg_in.rd_val.v = s.renamed_.rd_val
  //         # Copy over the non-opaque fields
  //         s.iq_slot_in.src0.v = s.renamed_.rs1
  //         s.iq_slot_in.src0_val.v = s.renamed_.rs1_val
  //         s.iq_slot_in.src1.v = s.renamed_.rs2
  //         s.iq_slot_in.src1_val.v = s.renamed_.rs2_val
  //         # Set the current readyness
  //         s.iq_slot_in.src0_rdy.v = s.is_ready_ready[0]
  //         s.iq_slot_in.src1_rdy.v = s.is_ready_ready[1]
  //
  //       s.iq.add_value.v = s.iq_slot_in
  //       s.iq.add_value.opaque.v = s.iq_msg_in

  // logic for handle_input()
  always @ (*) begin
    iq_slot_in = 0;
    iq_msg_in = 0;
    iq_msg_in[(74)-1:0] = renamed_[(74)-1:0];
    iq_slot_in[(2)-1:0] = renamed_[(74)-1:72];
    if ((renamed_[(2)-1:0] != PIPELINE_MSG_STATUS_VALID)) begin
      iq_slot_in[(160)-1:159] = 0;
      iq_slot_in[(152)-1:151] = 0;
      iq_msg_in[(142)-1:74] = renamed_[(142)-1:74];
    end
    else begin
      iq_msg_in[(135)-1:95] = renamed_[(135)-1:95];
      iq_msg_in[(95)-1:89] = renamed_[(95)-1:89];
      iq_msg_in[(89)-1:88] = renamed_[(89)-1:88];
      iq_slot_in[(158)-1:152] = renamed_[(81)-1:75];
      iq_slot_in[(160)-1:159] = renamed_[(75)-1:74];
      iq_slot_in[(150)-1:144] = renamed_[(88)-1:82];
      iq_slot_in[(152)-1:151] = renamed_[(82)-1:81];
      iq_slot_in[(159)-1:158] = is_ready_ready[0];
      iq_slot_in[(151)-1:150] = is_ready_ready[1];
    end
    iq$add_value = iq_slot_in;
    iq$add_value[(144)-1:2] = iq_msg_in;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_output():
  //       # Copy over the source info again
  //       s.peek_msg.v = 0
  //       s.peek_msg.v = s.iq.remove_value.opaque
  //       s.peek_msg.rs1.v = s.iq.remove_value.src0
  //       s.peek_msg.rs1_val.v = s.iq.remove_value.src0_val
  //       s.peek_msg.rs2.v = s.iq.remove_value.src1
  //       s.peek_msg.rs2_val.v = s.iq.remove_value.src1_val
  //       s.peek_msg.hdr_branch_mask.v = s.iq.remove_value.kill_opaque

  // logic for handle_output()
  always @ (*) begin
    peek_msg = 0;
    peek_msg = iq$remove_value[(144)-1:2];
    peek_msg[(81)-1:75] = iq$remove_value[(158)-1:152];
    peek_msg[(75)-1:74] = iq$remove_value[(160)-1:159];
    peek_msg[(88)-1:82] = iq$remove_value[(150)-1:144];
    peek_msg[(82)-1:81] = iq$remove_value[(152)-1:151];
    peek_msg[(74)-1:72] = iq$remove_value[(2)-1:0];
  end


endmodule // Issue_0x52678fcc1604a432

//-----------------------------------------------------------------------------
// CompactingIssueQueue_0x3a43583a53afd5b2
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.issue_queue {"interface": "add <CR> (value: Bits(160)) -> (); remove <CR> () -> (value: Bits(160)); notify <C> (value: Bits(6)) -> (); kill_notify (msg: Bits(5)) -> ()", "make_kill": "<function make_kill at 0x7f0068e319b0>", "num_slots": 2}
// PyMTL: verilator_xinit = zeros
module CompactingIssueQueue_0x3a43583a53afd5b2
(
  input  logic [   0:0] add_call,
  output logic  [   0:0] add_rdy,
  input  logic [ 159:0] add_value,
  input  logic [   0:0] clk,
  input  logic [   4:0] kill_notify_msg,
  input  logic [   0:0] notify_call,
  input  logic [   5:0] notify_value,
  input  logic [   0:0] remove_call,
  output logic  [   0:0] remove_rdy,
  output logic  [ 159:0] remove_value,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] do_shift_$000;
  logic   [   0:0] will_issue_$000;
  logic   [   0:0] will_issue_$001;


  // register declarations
  logic    [ 159:0] last_slot_in_;

  // localparam declarations
  localparam num_slots = 2;

  // loop variable declarations
  integer i;

  // slot_select_ temporaries
  logic   [   0:0] slot_select_$clk;
  logic   [   0:0] slot_select_$reset;
  logic   [   1:0] slot_select_$decode_signal;
  logic   [   0:0] slot_select_$decode_valid;
  logic   [   0:0] slot_select_$decode_decoded;

  PriorityDecoder_0x86563bd99c43c59 slot_select_
  (
    .clk            ( slot_select_$clk ),
    .reset          ( slot_select_$reset ),
    .decode_signal  ( slot_select_$decode_signal ),
    .decode_valid   ( slot_select_$decode_valid ),
    .decode_decoded ( slot_select_$decode_decoded )
  );

  // pdecode_packer_ temporaries
  logic   [   0:0] pdecode_packer_$clk;
  logic   [   0:0] pdecode_packer_$pack_in_$000;
  logic   [   0:0] pdecode_packer_$pack_in_$001;
  logic   [   0:0] pdecode_packer_$reset;
  logic   [   1:0] pdecode_packer_$pack_packed;

  Packer_0x67209f7520cf166 pdecode_packer_
  (
    .clk          ( pdecode_packer_$clk ),
    .pack_in_$000 ( pdecode_packer_$pack_in_$000 ),
    .pack_in_$001 ( pdecode_packer_$pack_in_$001 ),
    .reset        ( pdecode_packer_$reset ),
    .pack_packed  ( pdecode_packer_$pack_packed )
  );

  // slots_$000 temporaries
  logic   [ 159:0] slots_$000$input_value;
  logic   [   0:0] slots_$000$output_call;
  logic   [   0:0] slots_$000$clk;
  logic   [   4:0] slots_$000$kill_notify_msg;
  logic   [   5:0] slots_$000$notify_value;
  logic   [   0:0] slots_$000$input_call;
  logic   [   0:0] slots_$000$reset;
  logic   [   0:0] slots_$000$notify_call;
  logic   [   0:0] slots_$000$valid_ret;
  logic   [ 159:0] slots_$000$output_value;
  logic   [   0:0] slots_$000$ready_ret;

  GenericIssueSlot_0x3922269b2b56c3c3 slots_$000
  (
    .input_value     ( slots_$000$input_value ),
    .output_call     ( slots_$000$output_call ),
    .clk             ( slots_$000$clk ),
    .kill_notify_msg ( slots_$000$kill_notify_msg ),
    .notify_value    ( slots_$000$notify_value ),
    .input_call      ( slots_$000$input_call ),
    .reset           ( slots_$000$reset ),
    .notify_call     ( slots_$000$notify_call ),
    .valid_ret       ( slots_$000$valid_ret ),
    .output_value    ( slots_$000$output_value ),
    .ready_ret       ( slots_$000$ready_ret )
  );

  // slots_$001 temporaries
  logic   [ 159:0] slots_$001$input_value;
  logic   [   0:0] slots_$001$output_call;
  logic   [   0:0] slots_$001$clk;
  logic   [   4:0] slots_$001$kill_notify_msg;
  logic   [   5:0] slots_$001$notify_value;
  logic   [   0:0] slots_$001$input_call;
  logic   [   0:0] slots_$001$reset;
  logic   [   0:0] slots_$001$notify_call;
  logic   [   0:0] slots_$001$valid_ret;
  logic   [ 159:0] slots_$001$output_value;
  logic   [   0:0] slots_$001$ready_ret;

  GenericIssueSlot_0x3922269b2b56c3c3 slots_$001
  (
    .input_value     ( slots_$001$input_value ),
    .output_call     ( slots_$001$output_call ),
    .clk             ( slots_$001$clk ),
    .kill_notify_msg ( slots_$001$kill_notify_msg ),
    .notify_value    ( slots_$001$notify_value ),
    .input_call      ( slots_$001$input_call ),
    .reset           ( slots_$001$reset ),
    .notify_call     ( slots_$001$notify_call ),
    .valid_ret       ( slots_$001$valid_ret ),
    .output_value    ( slots_$001$output_value ),
    .ready_ret       ( slots_$001$ready_ret )
  );

  // mux_ temporaries
  logic   [ 159:0] mux_$mux_in_$000;
  logic   [ 159:0] mux_$mux_in_$001;
  logic   [   0:0] mux_$clk;
  logic   [   0:0] mux_$reset;
  logic   [   0:0] mux_$mux_select;
  logic   [ 159:0] mux_$mux_out;

  Mux_0x554c2b8bcd5014d5 mux_
  (
    .mux_in_$000 ( mux_$mux_in_$000 ),
    .mux_in_$001 ( mux_$mux_in_$001 ),
    .clk         ( mux_$clk ),
    .reset       ( mux_$reset ),
    .mux_select  ( mux_$mux_select ),
    .mux_out     ( mux_$mux_out )
  );

  // slot_issue_ temporaries
  logic   [   0:0] slot_issue_$clk;
  logic   [   0:0] slot_issue_$reset;
  logic   [   0:0] slot_issue_$encode_number;
  logic   [   1:0] slot_issue_$encode_onehot;

  OneHotEncoder_0x62af1c1ff9e32b51 slot_issue_
  (
    .clk           ( slot_issue_$clk ),
    .reset         ( slot_issue_$reset ),
    .encode_number ( slot_issue_$encode_number ),
    .encode_onehot ( slot_issue_$encode_onehot )
  );

  // signal connections
  assign mux_$clk                     = clk;
  assign mux_$mux_in_$000             = slots_$000$output_value;
  assign mux_$mux_in_$001             = slots_$001$output_value;
  assign mux_$mux_select              = slot_select_$decode_decoded;
  assign mux_$reset                   = reset;
  assign pdecode_packer_$clk          = clk;
  assign pdecode_packer_$pack_in_$000 = slots_$000$ready_ret;
  assign pdecode_packer_$pack_in_$001 = slots_$001$ready_ret;
  assign pdecode_packer_$reset        = reset;
  assign slot_issue_$clk              = clk;
  assign slot_issue_$encode_number    = slot_select_$decode_decoded;
  assign slot_issue_$reset            = reset;
  assign slot_select_$clk             = clk;
  assign slot_select_$decode_signal   = pdecode_packer_$pack_packed;
  assign slot_select_$decode_signal   = pdecode_packer_$pack_packed;
  assign slot_select_$reset           = reset;
  assign slots_$000$clk               = clk;
  assign slots_$000$kill_notify_msg   = kill_notify_msg;
  assign slots_$000$notify_call       = notify_call;
  assign slots_$000$notify_value      = notify_value;
  assign slots_$000$reset             = reset;
  assign slots_$001$clk               = clk;
  assign slots_$001$kill_notify_msg   = kill_notify_msg;
  assign slots_$001$notify_call       = notify_call;
  assign slots_$001$notify_value      = notify_value;
  assign slots_$001$reset             = reset;

  // array declarations
  logic    [   0:0] do_shift_[0:0];
  assign do_shift_$000 = do_shift_[  0];
  logic    [   0:0] slots_$input_call[0:1];
  assign slots_$000$input_call = slots_$input_call[  0];
  assign slots_$001$input_call = slots_$input_call[  1];
  logic    [ 159:0] slots_$input_value[0:1];
  assign slots_$000$input_value = slots_$input_value[  0];
  assign slots_$001$input_value = slots_$input_value[  1];
  logic    [   0:0] slots_$output_call[0:1];
  assign slots_$000$output_call = slots_$output_call[  0];
  assign slots_$001$output_call = slots_$output_call[  1];
  logic   [ 159:0] slots_$output_value[0:1];
  assign slots_$output_value[  0] = slots_$000$output_value;
  assign slots_$output_value[  1] = slots_$001$output_value;
  logic   [   0:0] slots_$valid_ret[0:1];
  assign slots_$valid_ret[  0] = slots_$000$valid_ret;
  assign slots_$valid_ret[  1] = slots_$001$valid_ret;
  logic    [   0:0] will_issue_[0:1];
  assign will_issue_$000 = will_issue_[  0];
  assign will_issue_$001 = will_issue_[  1];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def last_slot_input():
  //       s.slots_[num_slots - 1].input_value.v = s.last_slot_in_.v

  // logic for last_slot_input()
  always @ (*) begin
    slots_$input_value[(num_slots-1)] = last_slot_in_;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def slot_input(i=i):
  //         s.slots_[i].input_call.v = s.do_shift_[i]
  //         s.slots_[i].input_value.v = s.slots_[i + 1].output_value

  // logic for slot_input()
  always @ (*) begin
    slots_$input_call[0] = do_shift_[0];
    slots_$input_value[0] = slots_$output_value[(0+1)];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_add():
  //       # TODO: The kills from this cycle need to be forwarded to this:
  //       s.slots_[num_slots - 1].input_call.v = s.add_call
  //       s.last_slot_in_.v = s.add_value
  //       # Forward any notifications from current cycle
  //       if s.notify_call:
  //         if s.notify_value == s.add_value.src0:
  //           s.last_slot_in_.src0_rdy.v = 1
  //         if s.notify_value == s.add_value.src1:
  //           s.last_slot_in_.src1_rdy.v = 1

  // logic for handle_add()
  always @ (*) begin
    slots_$input_call[(num_slots-1)] = add_call;
    last_slot_in_ = add_value;
    if (notify_call) begin
      if ((notify_value == add_value[(158)-1:152])) begin
        last_slot_in_[(159)-1:158] = 1;
      end
      else begin
      end
      if ((notify_value == add_value[(150)-1:144])) begin
        last_slot_in_[(151)-1:150] = 1;
      end
      else begin
      end
    end
    else begin
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def shift0():
  //         # The 0th slot only shifts in if invalid or issuing
  //         s.do_shift_[0].v = (not s.slots_[0].valid_ret or
  //                             s.will_issue_[0]) and (s.slots_[1].valid_ret and
  //                                                    not s.will_issue_[1])

  // logic for shift0()
  always @ (*) begin
    do_shift_[0] = ((!slots_$valid_ret[0]||will_issue_[0])&&(slots_$valid_ret[1]&&!will_issue_[1]));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def output0():
  //       # The 0th slot only outputs if issuing
  //       s.slots_[0].output_call.v = s.will_issue_[0]

  // logic for output0()
  always @ (*) begin
    slots_$output_call[0] = will_issue_[0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def outputk(i=i):
  //         s.slots_[i].output_call.v = s.will_issue_[i] or s.do_shift_[i - 1]

  // logic for outputk()
  always @ (*) begin
    slots_$output_call[1] = (will_issue_[1]||do_shift_[(1-1)]);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def add_rdy():
  //       s.add_rdy.v = not s.slots_[num_slots - 1].valid_ret or s.slots_[
  //           num_slots - 1].output_call

  // logic for add_rdy()
  always @ (*) begin
    add_rdy = (!slots_$valid_ret[(num_slots-1)]||slots_$output_call[(num_slots-1)]);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_remove():
  //       s.remove_rdy.v = s.slot_select_.decode_valid
  //       s.remove_value.v = s.mux_.mux_out
  //       for i in range(num_slots):
  //         s.will_issue_[i].v = (
  //             s.slot_select_.decode_valid and s.remove_call and
  //             s.slot_issue_.encode_onehot[i])

  // logic for handle_remove()
  always @ (*) begin
    remove_rdy = slot_select_$decode_valid;
    remove_value = mux_$mux_out;
    for (i=0; i < num_slots; i=i+1)
    begin
      will_issue_[i] = (slot_select_$decode_valid&&remove_call&&slot_issue_$encode_onehot[i]);
    end
  end


endmodule // CompactingIssueQueue_0x3a43583a53afd5b2

//-----------------------------------------------------------------------------
// PriorityDecoder_0x86563bd99c43c59
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.coders {"inwidth": 2}
// PyMTL: verilator_xinit = zeros
module PriorityDecoder_0x86563bd99c43c59
(
  input  logic [   0:0] clk,
  output logic [   0:0] decode_decoded,
  input  logic [   1:0] decode_signal,
  output logic [   0:0] decode_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] outs$000;
  logic   [   0:0] outs$001;
  logic   [   0:0] outs$002;
  logic   [   0:0] valid$000;
  logic   [   0:0] valid$001;
  logic   [   0:0] valid$002;


  // signal connections
  assign decode_decoded = outs$002;
  assign decode_valid   = valid$002;
  assign outs$000       = 1'd0;
  assign valid$000      = 1'd0;

  // array declarations
  logic    [   0:0] outs[0:2];
  assign outs$000 = outs[  0];
  assign outs$001 = outs[  1];
  assign outs$002 = outs[  2];
  logic    [   0:0] valid[0:2];
  assign valid$000 = valid[  0];
  assign valid$001 = valid[  1];
  assign valid$002 = valid[  2];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[0]) begin
      valid[1] = 1;
      outs[1] = outs[0];
    end
    else begin
      if (decode_signal[0]) begin
        valid[1] = 1;
        outs[1] = 0;
      end
      else begin
        valid[1] = 0;
        outs[1] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[1]) begin
      valid[2] = 1;
      outs[2] = outs[1];
    end
    else begin
      if (decode_signal[1]) begin
        valid[2] = 1;
        outs[2] = 1;
      end
      else begin
        valid[2] = 0;
        outs[2] = 0;
      end
    end
  end


endmodule // PriorityDecoder_0x86563bd99c43c59

//-----------------------------------------------------------------------------
// Packer_0x67209f7520cf166
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.packers {"dtype": 1, "nports": 2}
// PyMTL: verilator_xinit = zeros
module Packer_0x67209f7520cf166
(
  input  logic [   0:0] clk,
  input  logic [   0:0] pack_in_$000,
  input  logic [   0:0] pack_in_$001,
  output logic  [   1:0] pack_packed,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nbits = 1;


  // array declarations
  logic   [   0:0] pack_in_[0:1];
  assign pack_in_[  0] = pack_in_$000;
  assign pack_in_[  1] = pack_in_$001;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(1)-1:0] = pack_in_[0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(2)-1:1] = pack_in_[1];
  end


endmodule // Packer_0x67209f7520cf166

//-----------------------------------------------------------------------------
// GenericIssueSlot_0x3922269b2b56c3c3
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.issue_queue {"interface": "kill_notify (msg: Bits(5)) -> (); notify <C> (value: Bits(6)) -> (); valid () -> (ret: Bits(1)); ready () -> (ret: Bits(1)); output <C> () -> (value: Bits(160)); input <C> (value: Bits(160)) -> ()", "make_kill": "<function make_kill at 0x7f0068e319b0>"}
// PyMTL: verilator_xinit = zeros
module GenericIssueSlot_0x3922269b2b56c3c3
(
  input  logic [   0:0] clk,
  input  logic [   0:0] input_call,
  input  logic [ 159:0] input_value,
  input  logic [   4:0] kill_notify_msg,
  input  logic [   0:0] notify_call,
  input  logic [   5:0] notify_value,
  input  logic [   0:0] output_call,
  output logic  [ 159:0] output_value,
  output logic  [   0:0] ready_ret,
  input  logic [   0:0] reset,
  output logic [   0:0] valid_ret
);

  // logic declarations
  logic   [   0:0] kill_;


  // register declarations
  logic    [   0:0] src0_match_;
  logic    [   0:0] src0_rdy_$write_call;
  logic    [   0:0] src0_rdy_$write_data;
  logic    [   0:0] src1_match_;
  logic    [   0:0] src1_rdy_$write_call;
  logic    [   0:0] src1_rdy_$write_data;
  logic    [   0:0] srcs_ready_;

  // src0_rdy_ temporaries
  logic   [   0:0] src0_rdy_$clk;
  logic   [   0:0] src0_rdy_$reset;
  logic   [   0:0] src0_rdy_$read_data;

  Register_0x6d252b2adb6c8882 src0_rdy_
  (
    .clk        ( src0_rdy_$clk ),
    .write_call ( src0_rdy_$write_call ),
    .write_data ( src0_rdy_$write_data ),
    .reset      ( src0_rdy_$reset ),
    .read_data  ( src0_rdy_$read_data )
  );

  // src1_val_ temporaries
  logic   [   0:0] src1_val_$clk;
  logic   [   0:0] src1_val_$write_call;
  logic   [   0:0] src1_val_$write_data;
  logic   [   0:0] src1_val_$reset;
  logic   [   0:0] src1_val_$read_data;

  Register_0x6d252b2adb6c8882 src1_val_
  (
    .clk        ( src1_val_$clk ),
    .write_call ( src1_val_$write_call ),
    .write_data ( src1_val_$write_data ),
    .reset      ( src1_val_$reset ),
    .read_data  ( src1_val_$read_data )
  );

  // src0_ temporaries
  logic   [   0:0] src0_$clk;
  logic   [   0:0] src0_$write_call;
  logic   [   5:0] src0_$write_data;
  logic   [   0:0] src0_$reset;
  logic   [   5:0] src0_$read_data;

  Register_0x44ce0714c41c17d4 src0_
  (
    .clk        ( src0_$clk ),
    .write_call ( src0_$write_call ),
    .write_data ( src0_$write_data ),
    .reset      ( src0_$reset ),
    .read_data  ( src0_$read_data )
  );

  // src1_rdy_ temporaries
  logic   [   0:0] src1_rdy_$clk;
  logic   [   0:0] src1_rdy_$reset;
  logic   [   0:0] src1_rdy_$read_data;

  Register_0x6d252b2adb6c8882 src1_rdy_
  (
    .clk        ( src1_rdy_$clk ),
    .write_call ( src1_rdy_$write_call ),
    .write_data ( src1_rdy_$write_data ),
    .reset      ( src1_rdy_$reset ),
    .read_data  ( src1_rdy_$read_data )
  );

  // val_manager_ temporaries
  logic   [   4:0] val_manager_$kill_notify_msg;
  logic   [   0:0] val_manager_$clk;
  logic   [   1:0] val_manager_$add_msg;
  logic   [   0:0] val_manager_$reset;
  logic   [   0:0] val_manager_$add_call;
  logic   [   0:0] val_manager_$take_call;
  logic   [   1:0] val_manager_$peek_msg;
  logic   [   0:0] val_manager_$add_rdy;
  logic   [   0:0] val_manager_$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb val_manager_
  (
    .kill_notify_msg ( val_manager_$kill_notify_msg ),
    .clk             ( val_manager_$clk ),
    .add_msg         ( val_manager_$add_msg ),
    .reset           ( val_manager_$reset ),
    .add_call        ( val_manager_$add_call ),
    .take_call       ( val_manager_$take_call ),
    .peek_msg        ( val_manager_$peek_msg ),
    .add_rdy         ( val_manager_$add_rdy ),
    .peek_rdy        ( val_manager_$peek_rdy )
  );

  // src1_ temporaries
  logic   [   0:0] src1_$clk;
  logic   [   0:0] src1_$write_call;
  logic   [   5:0] src1_$write_data;
  logic   [   0:0] src1_$reset;
  logic   [   5:0] src1_$read_data;

  Register_0x44ce0714c41c17d4 src1_
  (
    .clk        ( src1_$clk ),
    .write_call ( src1_$write_call ),
    .write_data ( src1_$write_data ),
    .reset      ( src1_$reset ),
    .read_data  ( src1_$read_data )
  );

  // src0_val_ temporaries
  logic   [   0:0] src0_val_$clk;
  logic   [   0:0] src0_val_$write_call;
  logic   [   0:0] src0_val_$write_data;
  logic   [   0:0] src0_val_$reset;
  logic   [   0:0] src0_val_$read_data;

  Register_0x6d252b2adb6c8882 src0_val_
  (
    .clk        ( src0_val_$clk ),
    .write_call ( src0_val_$write_call ),
    .write_data ( src0_val_$write_data ),
    .reset      ( src0_val_$reset ),
    .read_data  ( src0_val_$read_data )
  );

  // opaque_ temporaries
  logic   [   0:0] opaque_$clk;
  logic   [   0:0] opaque_$write_call;
  logic   [ 141:0] opaque_$write_data;
  logic   [   0:0] opaque_$reset;
  logic   [ 141:0] opaque_$read_data;

  Register_0x24d6bb878320116e opaque_
  (
    .clk        ( opaque_$clk ),
    .write_call ( opaque_$write_call ),
    .write_data ( opaque_$write_data ),
    .reset      ( opaque_$reset ),
    .read_data  ( opaque_$read_data )
  );

  // signal connections
  assign opaque_$clk                  = clk;
  assign opaque_$reset                = reset;
  assign opaque_$write_call           = input_call;
  assign opaque_$write_data           = input_value[143:2];
  assign output_value[143:2]          = opaque_$read_data;
  assign output_value[149:144]        = src1_$read_data;
  assign output_value[151:151]        = src1_val_$read_data;
  assign output_value[157:152]        = src0_$read_data;
  assign output_value[159:159]        = src0_val_$read_data;
  assign output_value[1:0]            = val_manager_$peek_msg;
  assign src0_$clk                    = clk;
  assign src0_$reset                  = reset;
  assign src0_$write_call             = input_call;
  assign src0_$write_data             = input_value[157:152];
  assign src0_rdy_$clk                = clk;
  assign src0_rdy_$reset              = reset;
  assign src0_val_$clk                = clk;
  assign src0_val_$reset              = reset;
  assign src0_val_$write_call         = input_call;
  assign src0_val_$write_data         = input_value[159:159];
  assign src1_$clk                    = clk;
  assign src1_$reset                  = reset;
  assign src1_$write_call             = input_call;
  assign src1_$write_data             = input_value[149:144];
  assign src1_rdy_$clk                = clk;
  assign src1_rdy_$reset              = reset;
  assign src1_val_$clk                = clk;
  assign src1_val_$reset              = reset;
  assign src1_val_$write_call         = input_call;
  assign src1_val_$write_data         = input_value[151:151];
  assign val_manager_$add_call        = input_call;
  assign val_manager_$add_msg         = input_value[1:0];
  assign val_manager_$clk             = clk;
  assign val_manager_$kill_notify_msg = kill_notify_msg;
  assign val_manager_$reset           = reset;
  assign val_manager_$take_call       = output_call;
  assign valid_ret                    = val_manager_$peek_rdy;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def match_src():
  //       s.src0_match_.v = s.src0_val_.read_data and s.notify_call and (
  //           s.src0_.read_data == s.notify_value)
  //       s.src1_match_.v = s.src1_val_.read_data and s.notify_call and (
  //           s.src1_.read_data == s.notify_value)

  // logic for match_src()
  always @ (*) begin
    src0_match_ = (src0_val_$read_data&&notify_call&&(src0_$read_data == notify_value));
    src1_match_ = (src1_val_$read_data&&notify_call&&(src1_$read_data == notify_value));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_outputs():
  //       s.output_value.src0_rdy.v = s.src0_rdy_.read_data or s.src0_match_
  //       s.output_value.src1_rdy.v = s.src1_rdy_.read_data or s.src1_match_
  //       s.srcs_ready_.v = s.output_value.src0_rdy and s.output_value.src1_rdy
  //       s.ready_ret.v = s.valid_ret and s.srcs_ready_

  // logic for handle_outputs()
  always @ (*) begin
    output_value[(159)-1:158] = (src0_rdy_$read_data||src0_match_);
    output_value[(151)-1:150] = (src1_rdy_$read_data||src1_match_);
    srcs_ready_ = (output_value[(159)-1:158]&&output_value[(151)-1:150]);
    ready_ret = (valid_ret&&srcs_ready_);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_rdy():
  //       s.src0_rdy_.write_call.v = s.input_call or (s.src0_match_ and s.valid_ret)
  //       s.src1_rdy_.write_call.v = s.input_call or (s.src1_match_ and s.valid_ret)
  //
  //       if s.input_call:
  //         s.src0_rdy_.write_data.v = s.input_value.src0_rdy or not s.input_value.src0_val
  //         s.src1_rdy_.write_data.v = s.input_value.src1_rdy or not s.input_value.src1_val
  //       else:
  //         s.src0_rdy_.write_data.v = s.src0_match_
  //         s.src1_rdy_.write_data.v = s.src1_match_

  // logic for set_rdy()
  always @ (*) begin
    src0_rdy_$write_call = (input_call||(src0_match_&&valid_ret));
    src1_rdy_$write_call = (input_call||(src1_match_&&valid_ret));
    if (input_call) begin
      src0_rdy_$write_data = (input_value[(159)-1:158]||!input_value[(160)-1:159]);
      src1_rdy_$write_data = (input_value[(151)-1:150]||!input_value[(152)-1:151]);
    end
    else begin
      src0_rdy_$write_data = src0_match_;
      src1_rdy_$write_data = src1_match_;
    end
  end


endmodule // GenericIssueSlot_0x3922269b2b56c3c3

//-----------------------------------------------------------------------------
// Register_0x6d252b2adb6c8882
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(1)); write <C> (data: Bits(1)) -> ()", "reset_value": null}
// PyMTL: verilator_xinit = zeros
module Register_0x6d252b2adb6c8882
(
  input  logic [   0:0] clk,
  output logic [   0:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [   0:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [   0:0] reg_value;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (update) begin
      reg_value <= write_data;
    end
    else begin
    end
  end


endmodule // Register_0x6d252b2adb6c8882

//-----------------------------------------------------------------------------
// Register_0x44ce0714c41c17d4
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(6)); write <C> (data: Bits(6)) -> ()", "reset_value": null}
// PyMTL: verilator_xinit = zeros
module Register_0x44ce0714c41c17d4
(
  input  logic [   0:0] clk,
  output logic [   5:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [   5:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [   5:0] reg_value;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (update) begin
      reg_value <= write_data;
    end
    else begin
    end
  end


endmodule // Register_0x44ce0714c41c17d4

//-----------------------------------------------------------------------------
// GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {}
// PyMTL: verilator_xinit = zeros
module GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb
(
  input  logic [   0:0] add_call,
  input  logic [   1:0] add_msg,
  output logic [   0:0] add_rdy,
  input  logic [   0:0] clk,
  input  logic [   4:0] kill_notify_msg,
  output logic [   1:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // manager temporaries
  logic   [   0:0] manager$check_keep;
  logic   [   0:0] manager$clk;
  logic   [   4:0] manager$kill_notify_msg;
  logic   [   1:0] manager$add_msg;
  logic   [   1:0] manager$check_out;
  logic   [   0:0] manager$reset;
  logic   [   0:0] manager$add_call;
  logic   [   0:0] manager$take_call;
  logic   [   1:0] manager$check_in_;
  logic   [   1:0] manager$peek_msg;
  logic   [   0:0] manager$add_rdy;
  logic   [   4:0] manager$check_msg;
  logic   [   0:0] manager$peek_rdy;

  ValidValueManager_0x335daa45f6084ab9 manager
  (
    .check_keep      ( manager$check_keep ),
    .clk             ( manager$clk ),
    .kill_notify_msg ( manager$kill_notify_msg ),
    .add_msg         ( manager$add_msg ),
    .check_out       ( manager$check_out ),
    .reset           ( manager$reset ),
    .add_call        ( manager$add_call ),
    .take_call       ( manager$take_call ),
    .check_in_       ( manager$check_in_ ),
    .peek_msg        ( manager$peek_msg ),
    .add_rdy         ( manager$add_rdy ),
    .check_msg       ( manager$check_msg ),
    .peek_rdy        ( manager$peek_rdy )
  );

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [   1:0] drop_controller$check_in_;
  logic   [   4:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [   1:0] drop_controller$check_out;

  KillDropController_0xccf15b584e8c1d drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // signal connections
  assign add_rdy                   = manager$add_rdy;
  assign drop_controller$check_in_ = manager$check_in_;
  assign drop_controller$check_msg = manager$check_msg;
  assign drop_controller$clk       = clk;
  assign drop_controller$reset     = reset;
  assign manager$add_call          = add_call;
  assign manager$add_msg           = add_msg;
  assign manager$check_keep        = drop_controller$check_keep;
  assign manager$check_out         = drop_controller$check_out;
  assign manager$clk               = clk;
  assign manager$kill_notify_msg   = kill_notify_msg;
  assign manager$reset             = reset;
  assign manager$take_call         = take_call;
  assign peek_msg                  = manager$peek_msg;
  assign peek_rdy                  = manager$peek_rdy;



endmodule // GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb

//-----------------------------------------------------------------------------
// ValidValueManager_0x335daa45f6084ab9
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"interface": "kill_notify (msg: Bits(5)) -> (); peek <R> () -> (msg: Bits(2)); take <C> () -> (); add <CR> (msg: Bits(2)) -> ()"}
// PyMTL: verilator_xinit = zeros
module ValidValueManager_0x335daa45f6084ab9
(
  input  logic [   0:0] add_call,
  input  logic [   1:0] add_msg,
  output logic [   0:0] add_rdy,
  output logic [   1:0] check_in_,
  input  logic [   0:0] check_keep,
  output logic [   4:0] check_msg,
  input  logic [   1:0] check_out,
  input  logic [   0:0] clk,
  input  logic [   4:0] kill_notify_msg,
  output logic [   1:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // register declarations
  logic    [   0:0] output_clear;
  logic    [   0:0] output_rdy;
  logic    [   0:0] val_reg$write_data;

  // val_reg temporaries
  logic   [   0:0] val_reg$clk;
  logic   [   0:0] val_reg$reset;
  logic   [   0:0] val_reg$read_data;

  Register_0x360ff20b8ea9d7d7 val_reg
  (
    .clk        ( val_reg$clk ),
    .write_data ( val_reg$write_data ),
    .reset      ( val_reg$reset ),
    .read_data  ( val_reg$read_data )
  );

  // out_reg temporaries
  logic   [   0:0] out_reg$clk;
  logic   [   0:0] out_reg$write_call;
  logic   [   1:0] out_reg$write_data;
  logic   [   0:0] out_reg$reset;
  logic   [   1:0] out_reg$read_data;

  Register_0x2ae482f34ea2364c out_reg
  (
    .clk        ( out_reg$clk ),
    .write_call ( out_reg$write_call ),
    .write_data ( out_reg$write_data ),
    .reset      ( out_reg$reset ),
    .read_data  ( out_reg$read_data )
  );

  // signal connections
  assign add_rdy            = output_clear;
  assign check_in_          = out_reg$read_data;
  assign check_msg          = kill_notify_msg;
  assign out_reg$clk        = clk;
  assign out_reg$reset      = reset;
  assign out_reg$write_call = add_call;
  assign out_reg$write_data = add_msg;
  assign peek_msg           = check_out;
  assign peek_rdy           = output_rdy;
  assign val_reg$clk        = clk;
  assign val_reg$reset      = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_rdy():
  //       if s.val_reg.read_data:
  //         s.output_rdy.v = s.check_keep
  //       else:
  //         s.output_rdy.v = 0

  // logic for handle_rdy()
  always @ (*) begin
    if (val_reg$read_data) begin
      output_rdy = check_keep;
    end
    else begin
      output_rdy = 0;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_clear():
  //       s.output_clear.v = not s.output_rdy or s.take_call

  // logic for handle_clear()
  always @ (*) begin
    output_clear = (!output_rdy||take_call);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_val_reg_in():
  //       if s.add_call:
  //         s.val_reg.write_data.v = 1
  //       else:
  //         s.val_reg.write_data.v = not s.output_clear

  // logic for handle_val_reg_in()
  always @ (*) begin
    if (add_call) begin
      val_reg$write_data = 1;
    end
    else begin
      val_reg$write_data = !output_clear;
    end
  end


endmodule // ValidValueManager_0x335daa45f6084ab9

//-----------------------------------------------------------------------------
// Register_0x2ae482f34ea2364c
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(2)); write <C> (data: Bits(2)) -> ()", "reset_value": null}
// PyMTL: verilator_xinit = zeros
module Register_0x2ae482f34ea2364c
(
  input  logic [   0:0] clk,
  output logic [   1:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [   1:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [   1:0] reg_value;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (update) begin
      reg_value <= write_data;
    end
    else begin
    end
  end


endmodule // Register_0x2ae482f34ea2364c

//-----------------------------------------------------------------------------
// Mux_0x554c2b8bcd5014d5
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.mux {"dtype": 160, "nports": 2}
// PyMTL: verilator_xinit = zeros
module Mux_0x554c2b8bcd5014d5
(
  input  logic [   0:0] clk,
  input  logic [ 159:0] mux_in_$000,
  input  logic [ 159:0] mux_in_$001,
  output logic  [ 159:0] mux_out,
  input  logic [   0:0] mux_select,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nports = 2;


  // array declarations
  logic   [ 159:0] mux_in_[0:1];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def select():
  //       assert s.mux_select < nports
  //       s.mux_out.v = s.mux_in_[s.mux_select]

  // logic for select()
  always @ (*) begin
    mux_out = mux_in_[mux_select];
  end


endmodule // Mux_0x554c2b8bcd5014d5

//-----------------------------------------------------------------------------
// OneHotEncoder_0x62af1c1ff9e32b51
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.onehot {"enable": false, "noutbits": 2}
// PyMTL: verilator_xinit = zeros
module OneHotEncoder_0x62af1c1ff9e32b51
(
  input  logic [   0:0] clk,
  input  logic [   0:0] encode_number,
  output logic  [   1:0] encode_onehot,
  input  logic [   0:0] reset
);



  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[0] = (encode_number == 0);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[1] = (encode_number == 1);
  end


endmodule // OneHotEncoder_0x62af1c1ff9e32b51

//-----------------------------------------------------------------------------
// PriorityDecoder_0x2e5c0266b409153a
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.coders {"inwidth": 64}
// PyMTL: verilator_xinit = zeros
module PriorityDecoder_0x2e5c0266b409153a
(
  input  logic [   0:0] clk,
  output logic [   5:0] decode_decoded,
  input  logic [  63:0] decode_signal,
  output logic [   0:0] decode_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   5:0] outs$000;
  logic   [   5:0] outs$001;
  logic   [   5:0] outs$002;
  logic   [   5:0] outs$003;
  logic   [   5:0] outs$004;
  logic   [   5:0] outs$005;
  logic   [   5:0] outs$006;
  logic   [   5:0] outs$007;
  logic   [   5:0] outs$008;
  logic   [   5:0] outs$009;
  logic   [   5:0] outs$010;
  logic   [   5:0] outs$011;
  logic   [   5:0] outs$012;
  logic   [   5:0] outs$013;
  logic   [   5:0] outs$014;
  logic   [   5:0] outs$015;
  logic   [   5:0] outs$016;
  logic   [   5:0] outs$017;
  logic   [   5:0] outs$018;
  logic   [   5:0] outs$019;
  logic   [   5:0] outs$020;
  logic   [   5:0] outs$021;
  logic   [   5:0] outs$022;
  logic   [   5:0] outs$023;
  logic   [   5:0] outs$024;
  logic   [   5:0] outs$025;
  logic   [   5:0] outs$026;
  logic   [   5:0] outs$027;
  logic   [   5:0] outs$028;
  logic   [   5:0] outs$029;
  logic   [   5:0] outs$030;
  logic   [   5:0] outs$031;
  logic   [   5:0] outs$032;
  logic   [   5:0] outs$033;
  logic   [   5:0] outs$034;
  logic   [   5:0] outs$035;
  logic   [   5:0] outs$036;
  logic   [   5:0] outs$037;
  logic   [   5:0] outs$038;
  logic   [   5:0] outs$039;
  logic   [   5:0] outs$040;
  logic   [   5:0] outs$041;
  logic   [   5:0] outs$042;
  logic   [   5:0] outs$043;
  logic   [   5:0] outs$044;
  logic   [   5:0] outs$045;
  logic   [   5:0] outs$046;
  logic   [   5:0] outs$047;
  logic   [   5:0] outs$048;
  logic   [   5:0] outs$049;
  logic   [   5:0] outs$050;
  logic   [   5:0] outs$051;
  logic   [   5:0] outs$052;
  logic   [   5:0] outs$053;
  logic   [   5:0] outs$054;
  logic   [   5:0] outs$055;
  logic   [   5:0] outs$056;
  logic   [   5:0] outs$057;
  logic   [   5:0] outs$058;
  logic   [   5:0] outs$059;
  logic   [   5:0] outs$060;
  logic   [   5:0] outs$061;
  logic   [   5:0] outs$062;
  logic   [   5:0] outs$063;
  logic   [   5:0] outs$064;
  logic   [   0:0] valid$000;
  logic   [   0:0] valid$001;
  logic   [   0:0] valid$002;
  logic   [   0:0] valid$003;
  logic   [   0:0] valid$004;
  logic   [   0:0] valid$005;
  logic   [   0:0] valid$006;
  logic   [   0:0] valid$007;
  logic   [   0:0] valid$008;
  logic   [   0:0] valid$009;
  logic   [   0:0] valid$010;
  logic   [   0:0] valid$011;
  logic   [   0:0] valid$012;
  logic   [   0:0] valid$013;
  logic   [   0:0] valid$014;
  logic   [   0:0] valid$015;
  logic   [   0:0] valid$016;
  logic   [   0:0] valid$017;
  logic   [   0:0] valid$018;
  logic   [   0:0] valid$019;
  logic   [   0:0] valid$020;
  logic   [   0:0] valid$021;
  logic   [   0:0] valid$022;
  logic   [   0:0] valid$023;
  logic   [   0:0] valid$024;
  logic   [   0:0] valid$025;
  logic   [   0:0] valid$026;
  logic   [   0:0] valid$027;
  logic   [   0:0] valid$028;
  logic   [   0:0] valid$029;
  logic   [   0:0] valid$030;
  logic   [   0:0] valid$031;
  logic   [   0:0] valid$032;
  logic   [   0:0] valid$033;
  logic   [   0:0] valid$034;
  logic   [   0:0] valid$035;
  logic   [   0:0] valid$036;
  logic   [   0:0] valid$037;
  logic   [   0:0] valid$038;
  logic   [   0:0] valid$039;
  logic   [   0:0] valid$040;
  logic   [   0:0] valid$041;
  logic   [   0:0] valid$042;
  logic   [   0:0] valid$043;
  logic   [   0:0] valid$044;
  logic   [   0:0] valid$045;
  logic   [   0:0] valid$046;
  logic   [   0:0] valid$047;
  logic   [   0:0] valid$048;
  logic   [   0:0] valid$049;
  logic   [   0:0] valid$050;
  logic   [   0:0] valid$051;
  logic   [   0:0] valid$052;
  logic   [   0:0] valid$053;
  logic   [   0:0] valid$054;
  logic   [   0:0] valid$055;
  logic   [   0:0] valid$056;
  logic   [   0:0] valid$057;
  logic   [   0:0] valid$058;
  logic   [   0:0] valid$059;
  logic   [   0:0] valid$060;
  logic   [   0:0] valid$061;
  logic   [   0:0] valid$062;
  logic   [   0:0] valid$063;
  logic   [   0:0] valid$064;


  // signal connections
  assign decode_decoded = outs$064;
  assign decode_valid   = valid$064;
  assign outs$000       = 6'd0;
  assign valid$000      = 1'd0;

  // array declarations
  logic    [   5:0] outs[0:64];
  assign outs$000 = outs[  0];
  assign outs$001 = outs[  1];
  assign outs$002 = outs[  2];
  assign outs$003 = outs[  3];
  assign outs$004 = outs[  4];
  assign outs$005 = outs[  5];
  assign outs$006 = outs[  6];
  assign outs$007 = outs[  7];
  assign outs$008 = outs[  8];
  assign outs$009 = outs[  9];
  assign outs$010 = outs[ 10];
  assign outs$011 = outs[ 11];
  assign outs$012 = outs[ 12];
  assign outs$013 = outs[ 13];
  assign outs$014 = outs[ 14];
  assign outs$015 = outs[ 15];
  assign outs$016 = outs[ 16];
  assign outs$017 = outs[ 17];
  assign outs$018 = outs[ 18];
  assign outs$019 = outs[ 19];
  assign outs$020 = outs[ 20];
  assign outs$021 = outs[ 21];
  assign outs$022 = outs[ 22];
  assign outs$023 = outs[ 23];
  assign outs$024 = outs[ 24];
  assign outs$025 = outs[ 25];
  assign outs$026 = outs[ 26];
  assign outs$027 = outs[ 27];
  assign outs$028 = outs[ 28];
  assign outs$029 = outs[ 29];
  assign outs$030 = outs[ 30];
  assign outs$031 = outs[ 31];
  assign outs$032 = outs[ 32];
  assign outs$033 = outs[ 33];
  assign outs$034 = outs[ 34];
  assign outs$035 = outs[ 35];
  assign outs$036 = outs[ 36];
  assign outs$037 = outs[ 37];
  assign outs$038 = outs[ 38];
  assign outs$039 = outs[ 39];
  assign outs$040 = outs[ 40];
  assign outs$041 = outs[ 41];
  assign outs$042 = outs[ 42];
  assign outs$043 = outs[ 43];
  assign outs$044 = outs[ 44];
  assign outs$045 = outs[ 45];
  assign outs$046 = outs[ 46];
  assign outs$047 = outs[ 47];
  assign outs$048 = outs[ 48];
  assign outs$049 = outs[ 49];
  assign outs$050 = outs[ 50];
  assign outs$051 = outs[ 51];
  assign outs$052 = outs[ 52];
  assign outs$053 = outs[ 53];
  assign outs$054 = outs[ 54];
  assign outs$055 = outs[ 55];
  assign outs$056 = outs[ 56];
  assign outs$057 = outs[ 57];
  assign outs$058 = outs[ 58];
  assign outs$059 = outs[ 59];
  assign outs$060 = outs[ 60];
  assign outs$061 = outs[ 61];
  assign outs$062 = outs[ 62];
  assign outs$063 = outs[ 63];
  assign outs$064 = outs[ 64];
  logic    [   0:0] valid[0:64];
  assign valid$000 = valid[  0];
  assign valid$001 = valid[  1];
  assign valid$002 = valid[  2];
  assign valid$003 = valid[  3];
  assign valid$004 = valid[  4];
  assign valid$005 = valid[  5];
  assign valid$006 = valid[  6];
  assign valid$007 = valid[  7];
  assign valid$008 = valid[  8];
  assign valid$009 = valid[  9];
  assign valid$010 = valid[ 10];
  assign valid$011 = valid[ 11];
  assign valid$012 = valid[ 12];
  assign valid$013 = valid[ 13];
  assign valid$014 = valid[ 14];
  assign valid$015 = valid[ 15];
  assign valid$016 = valid[ 16];
  assign valid$017 = valid[ 17];
  assign valid$018 = valid[ 18];
  assign valid$019 = valid[ 19];
  assign valid$020 = valid[ 20];
  assign valid$021 = valid[ 21];
  assign valid$022 = valid[ 22];
  assign valid$023 = valid[ 23];
  assign valid$024 = valid[ 24];
  assign valid$025 = valid[ 25];
  assign valid$026 = valid[ 26];
  assign valid$027 = valid[ 27];
  assign valid$028 = valid[ 28];
  assign valid$029 = valid[ 29];
  assign valid$030 = valid[ 30];
  assign valid$031 = valid[ 31];
  assign valid$032 = valid[ 32];
  assign valid$033 = valid[ 33];
  assign valid$034 = valid[ 34];
  assign valid$035 = valid[ 35];
  assign valid$036 = valid[ 36];
  assign valid$037 = valid[ 37];
  assign valid$038 = valid[ 38];
  assign valid$039 = valid[ 39];
  assign valid$040 = valid[ 40];
  assign valid$041 = valid[ 41];
  assign valid$042 = valid[ 42];
  assign valid$043 = valid[ 43];
  assign valid$044 = valid[ 44];
  assign valid$045 = valid[ 45];
  assign valid$046 = valid[ 46];
  assign valid$047 = valid[ 47];
  assign valid$048 = valid[ 48];
  assign valid$049 = valid[ 49];
  assign valid$050 = valid[ 50];
  assign valid$051 = valid[ 51];
  assign valid$052 = valid[ 52];
  assign valid$053 = valid[ 53];
  assign valid$054 = valid[ 54];
  assign valid$055 = valid[ 55];
  assign valid$056 = valid[ 56];
  assign valid$057 = valid[ 57];
  assign valid$058 = valid[ 58];
  assign valid$059 = valid[ 59];
  assign valid$060 = valid[ 60];
  assign valid$061 = valid[ 61];
  assign valid$062 = valid[ 62];
  assign valid$063 = valid[ 63];
  assign valid$064 = valid[ 64];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[0]) begin
      valid[1] = 1;
      outs[1] = outs[0];
    end
    else begin
      if (decode_signal[0]) begin
        valid[1] = 1;
        outs[1] = 0;
      end
      else begin
        valid[1] = 0;
        outs[1] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[1]) begin
      valid[2] = 1;
      outs[2] = outs[1];
    end
    else begin
      if (decode_signal[1]) begin
        valid[2] = 1;
        outs[2] = 1;
      end
      else begin
        valid[2] = 0;
        outs[2] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[2]) begin
      valid[3] = 1;
      outs[3] = outs[2];
    end
    else begin
      if (decode_signal[2]) begin
        valid[3] = 1;
        outs[3] = 2;
      end
      else begin
        valid[3] = 0;
        outs[3] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[3]) begin
      valid[4] = 1;
      outs[4] = outs[3];
    end
    else begin
      if (decode_signal[3]) begin
        valid[4] = 1;
        outs[4] = 3;
      end
      else begin
        valid[4] = 0;
        outs[4] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[4]) begin
      valid[5] = 1;
      outs[5] = outs[4];
    end
    else begin
      if (decode_signal[4]) begin
        valid[5] = 1;
        outs[5] = 4;
      end
      else begin
        valid[5] = 0;
        outs[5] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[5]) begin
      valid[6] = 1;
      outs[6] = outs[5];
    end
    else begin
      if (decode_signal[5]) begin
        valid[6] = 1;
        outs[6] = 5;
      end
      else begin
        valid[6] = 0;
        outs[6] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[6]) begin
      valid[7] = 1;
      outs[7] = outs[6];
    end
    else begin
      if (decode_signal[6]) begin
        valid[7] = 1;
        outs[7] = 6;
      end
      else begin
        valid[7] = 0;
        outs[7] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[7]) begin
      valid[8] = 1;
      outs[8] = outs[7];
    end
    else begin
      if (decode_signal[7]) begin
        valid[8] = 1;
        outs[8] = 7;
      end
      else begin
        valid[8] = 0;
        outs[8] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[8]) begin
      valid[9] = 1;
      outs[9] = outs[8];
    end
    else begin
      if (decode_signal[8]) begin
        valid[9] = 1;
        outs[9] = 8;
      end
      else begin
        valid[9] = 0;
        outs[9] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[9]) begin
      valid[10] = 1;
      outs[10] = outs[9];
    end
    else begin
      if (decode_signal[9]) begin
        valid[10] = 1;
        outs[10] = 9;
      end
      else begin
        valid[10] = 0;
        outs[10] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[10]) begin
      valid[11] = 1;
      outs[11] = outs[10];
    end
    else begin
      if (decode_signal[10]) begin
        valid[11] = 1;
        outs[11] = 10;
      end
      else begin
        valid[11] = 0;
        outs[11] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[11]) begin
      valid[12] = 1;
      outs[12] = outs[11];
    end
    else begin
      if (decode_signal[11]) begin
        valid[12] = 1;
        outs[12] = 11;
      end
      else begin
        valid[12] = 0;
        outs[12] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[12]) begin
      valid[13] = 1;
      outs[13] = outs[12];
    end
    else begin
      if (decode_signal[12]) begin
        valid[13] = 1;
        outs[13] = 12;
      end
      else begin
        valid[13] = 0;
        outs[13] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[13]) begin
      valid[14] = 1;
      outs[14] = outs[13];
    end
    else begin
      if (decode_signal[13]) begin
        valid[14] = 1;
        outs[14] = 13;
      end
      else begin
        valid[14] = 0;
        outs[14] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[14]) begin
      valid[15] = 1;
      outs[15] = outs[14];
    end
    else begin
      if (decode_signal[14]) begin
        valid[15] = 1;
        outs[15] = 14;
      end
      else begin
        valid[15] = 0;
        outs[15] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[15]) begin
      valid[16] = 1;
      outs[16] = outs[15];
    end
    else begin
      if (decode_signal[15]) begin
        valid[16] = 1;
        outs[16] = 15;
      end
      else begin
        valid[16] = 0;
        outs[16] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[16]) begin
      valid[17] = 1;
      outs[17] = outs[16];
    end
    else begin
      if (decode_signal[16]) begin
        valid[17] = 1;
        outs[17] = 16;
      end
      else begin
        valid[17] = 0;
        outs[17] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[17]) begin
      valid[18] = 1;
      outs[18] = outs[17];
    end
    else begin
      if (decode_signal[17]) begin
        valid[18] = 1;
        outs[18] = 17;
      end
      else begin
        valid[18] = 0;
        outs[18] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[18]) begin
      valid[19] = 1;
      outs[19] = outs[18];
    end
    else begin
      if (decode_signal[18]) begin
        valid[19] = 1;
        outs[19] = 18;
      end
      else begin
        valid[19] = 0;
        outs[19] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[19]) begin
      valid[20] = 1;
      outs[20] = outs[19];
    end
    else begin
      if (decode_signal[19]) begin
        valid[20] = 1;
        outs[20] = 19;
      end
      else begin
        valid[20] = 0;
        outs[20] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[20]) begin
      valid[21] = 1;
      outs[21] = outs[20];
    end
    else begin
      if (decode_signal[20]) begin
        valid[21] = 1;
        outs[21] = 20;
      end
      else begin
        valid[21] = 0;
        outs[21] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[21]) begin
      valid[22] = 1;
      outs[22] = outs[21];
    end
    else begin
      if (decode_signal[21]) begin
        valid[22] = 1;
        outs[22] = 21;
      end
      else begin
        valid[22] = 0;
        outs[22] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[22]) begin
      valid[23] = 1;
      outs[23] = outs[22];
    end
    else begin
      if (decode_signal[22]) begin
        valid[23] = 1;
        outs[23] = 22;
      end
      else begin
        valid[23] = 0;
        outs[23] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[23]) begin
      valid[24] = 1;
      outs[24] = outs[23];
    end
    else begin
      if (decode_signal[23]) begin
        valid[24] = 1;
        outs[24] = 23;
      end
      else begin
        valid[24] = 0;
        outs[24] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[24]) begin
      valid[25] = 1;
      outs[25] = outs[24];
    end
    else begin
      if (decode_signal[24]) begin
        valid[25] = 1;
        outs[25] = 24;
      end
      else begin
        valid[25] = 0;
        outs[25] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[25]) begin
      valid[26] = 1;
      outs[26] = outs[25];
    end
    else begin
      if (decode_signal[25]) begin
        valid[26] = 1;
        outs[26] = 25;
      end
      else begin
        valid[26] = 0;
        outs[26] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[26]) begin
      valid[27] = 1;
      outs[27] = outs[26];
    end
    else begin
      if (decode_signal[26]) begin
        valid[27] = 1;
        outs[27] = 26;
      end
      else begin
        valid[27] = 0;
        outs[27] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[27]) begin
      valid[28] = 1;
      outs[28] = outs[27];
    end
    else begin
      if (decode_signal[27]) begin
        valid[28] = 1;
        outs[28] = 27;
      end
      else begin
        valid[28] = 0;
        outs[28] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[28]) begin
      valid[29] = 1;
      outs[29] = outs[28];
    end
    else begin
      if (decode_signal[28]) begin
        valid[29] = 1;
        outs[29] = 28;
      end
      else begin
        valid[29] = 0;
        outs[29] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[29]) begin
      valid[30] = 1;
      outs[30] = outs[29];
    end
    else begin
      if (decode_signal[29]) begin
        valid[30] = 1;
        outs[30] = 29;
      end
      else begin
        valid[30] = 0;
        outs[30] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[30]) begin
      valid[31] = 1;
      outs[31] = outs[30];
    end
    else begin
      if (decode_signal[30]) begin
        valid[31] = 1;
        outs[31] = 30;
      end
      else begin
        valid[31] = 0;
        outs[31] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[31]) begin
      valid[32] = 1;
      outs[32] = outs[31];
    end
    else begin
      if (decode_signal[31]) begin
        valid[32] = 1;
        outs[32] = 31;
      end
      else begin
        valid[32] = 0;
        outs[32] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[32]) begin
      valid[33] = 1;
      outs[33] = outs[32];
    end
    else begin
      if (decode_signal[32]) begin
        valid[33] = 1;
        outs[33] = 32;
      end
      else begin
        valid[33] = 0;
        outs[33] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[33]) begin
      valid[34] = 1;
      outs[34] = outs[33];
    end
    else begin
      if (decode_signal[33]) begin
        valid[34] = 1;
        outs[34] = 33;
      end
      else begin
        valid[34] = 0;
        outs[34] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[34]) begin
      valid[35] = 1;
      outs[35] = outs[34];
    end
    else begin
      if (decode_signal[34]) begin
        valid[35] = 1;
        outs[35] = 34;
      end
      else begin
        valid[35] = 0;
        outs[35] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[35]) begin
      valid[36] = 1;
      outs[36] = outs[35];
    end
    else begin
      if (decode_signal[35]) begin
        valid[36] = 1;
        outs[36] = 35;
      end
      else begin
        valid[36] = 0;
        outs[36] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[36]) begin
      valid[37] = 1;
      outs[37] = outs[36];
    end
    else begin
      if (decode_signal[36]) begin
        valid[37] = 1;
        outs[37] = 36;
      end
      else begin
        valid[37] = 0;
        outs[37] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[37]) begin
      valid[38] = 1;
      outs[38] = outs[37];
    end
    else begin
      if (decode_signal[37]) begin
        valid[38] = 1;
        outs[38] = 37;
      end
      else begin
        valid[38] = 0;
        outs[38] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[38]) begin
      valid[39] = 1;
      outs[39] = outs[38];
    end
    else begin
      if (decode_signal[38]) begin
        valid[39] = 1;
        outs[39] = 38;
      end
      else begin
        valid[39] = 0;
        outs[39] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[39]) begin
      valid[40] = 1;
      outs[40] = outs[39];
    end
    else begin
      if (decode_signal[39]) begin
        valid[40] = 1;
        outs[40] = 39;
      end
      else begin
        valid[40] = 0;
        outs[40] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[40]) begin
      valid[41] = 1;
      outs[41] = outs[40];
    end
    else begin
      if (decode_signal[40]) begin
        valid[41] = 1;
        outs[41] = 40;
      end
      else begin
        valid[41] = 0;
        outs[41] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[41]) begin
      valid[42] = 1;
      outs[42] = outs[41];
    end
    else begin
      if (decode_signal[41]) begin
        valid[42] = 1;
        outs[42] = 41;
      end
      else begin
        valid[42] = 0;
        outs[42] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[42]) begin
      valid[43] = 1;
      outs[43] = outs[42];
    end
    else begin
      if (decode_signal[42]) begin
        valid[43] = 1;
        outs[43] = 42;
      end
      else begin
        valid[43] = 0;
        outs[43] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[43]) begin
      valid[44] = 1;
      outs[44] = outs[43];
    end
    else begin
      if (decode_signal[43]) begin
        valid[44] = 1;
        outs[44] = 43;
      end
      else begin
        valid[44] = 0;
        outs[44] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[44]) begin
      valid[45] = 1;
      outs[45] = outs[44];
    end
    else begin
      if (decode_signal[44]) begin
        valid[45] = 1;
        outs[45] = 44;
      end
      else begin
        valid[45] = 0;
        outs[45] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[45]) begin
      valid[46] = 1;
      outs[46] = outs[45];
    end
    else begin
      if (decode_signal[45]) begin
        valid[46] = 1;
        outs[46] = 45;
      end
      else begin
        valid[46] = 0;
        outs[46] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[46]) begin
      valid[47] = 1;
      outs[47] = outs[46];
    end
    else begin
      if (decode_signal[46]) begin
        valid[47] = 1;
        outs[47] = 46;
      end
      else begin
        valid[47] = 0;
        outs[47] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[47]) begin
      valid[48] = 1;
      outs[48] = outs[47];
    end
    else begin
      if (decode_signal[47]) begin
        valid[48] = 1;
        outs[48] = 47;
      end
      else begin
        valid[48] = 0;
        outs[48] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[48]) begin
      valid[49] = 1;
      outs[49] = outs[48];
    end
    else begin
      if (decode_signal[48]) begin
        valid[49] = 1;
        outs[49] = 48;
      end
      else begin
        valid[49] = 0;
        outs[49] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[49]) begin
      valid[50] = 1;
      outs[50] = outs[49];
    end
    else begin
      if (decode_signal[49]) begin
        valid[50] = 1;
        outs[50] = 49;
      end
      else begin
        valid[50] = 0;
        outs[50] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[50]) begin
      valid[51] = 1;
      outs[51] = outs[50];
    end
    else begin
      if (decode_signal[50]) begin
        valid[51] = 1;
        outs[51] = 50;
      end
      else begin
        valid[51] = 0;
        outs[51] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[51]) begin
      valid[52] = 1;
      outs[52] = outs[51];
    end
    else begin
      if (decode_signal[51]) begin
        valid[52] = 1;
        outs[52] = 51;
      end
      else begin
        valid[52] = 0;
        outs[52] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[52]) begin
      valid[53] = 1;
      outs[53] = outs[52];
    end
    else begin
      if (decode_signal[52]) begin
        valid[53] = 1;
        outs[53] = 52;
      end
      else begin
        valid[53] = 0;
        outs[53] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[53]) begin
      valid[54] = 1;
      outs[54] = outs[53];
    end
    else begin
      if (decode_signal[53]) begin
        valid[54] = 1;
        outs[54] = 53;
      end
      else begin
        valid[54] = 0;
        outs[54] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[54]) begin
      valid[55] = 1;
      outs[55] = outs[54];
    end
    else begin
      if (decode_signal[54]) begin
        valid[55] = 1;
        outs[55] = 54;
      end
      else begin
        valid[55] = 0;
        outs[55] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[55]) begin
      valid[56] = 1;
      outs[56] = outs[55];
    end
    else begin
      if (decode_signal[55]) begin
        valid[56] = 1;
        outs[56] = 55;
      end
      else begin
        valid[56] = 0;
        outs[56] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[56]) begin
      valid[57] = 1;
      outs[57] = outs[56];
    end
    else begin
      if (decode_signal[56]) begin
        valid[57] = 1;
        outs[57] = 56;
      end
      else begin
        valid[57] = 0;
        outs[57] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[57]) begin
      valid[58] = 1;
      outs[58] = outs[57];
    end
    else begin
      if (decode_signal[57]) begin
        valid[58] = 1;
        outs[58] = 57;
      end
      else begin
        valid[58] = 0;
        outs[58] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[58]) begin
      valid[59] = 1;
      outs[59] = outs[58];
    end
    else begin
      if (decode_signal[58]) begin
        valid[59] = 1;
        outs[59] = 58;
      end
      else begin
        valid[59] = 0;
        outs[59] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[59]) begin
      valid[60] = 1;
      outs[60] = outs[59];
    end
    else begin
      if (decode_signal[59]) begin
        valid[60] = 1;
        outs[60] = 59;
      end
      else begin
        valid[60] = 0;
        outs[60] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[60]) begin
      valid[61] = 1;
      outs[61] = outs[60];
    end
    else begin
      if (decode_signal[60]) begin
        valid[61] = 1;
        outs[61] = 60;
      end
      else begin
        valid[61] = 0;
        outs[61] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[61]) begin
      valid[62] = 1;
      outs[62] = outs[61];
    end
    else begin
      if (decode_signal[61]) begin
        valid[62] = 1;
        outs[62] = 61;
      end
      else begin
        valid[62] = 0;
        outs[62] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[62]) begin
      valid[63] = 1;
      outs[63] = outs[62];
    end
    else begin
      if (decode_signal[62]) begin
        valid[63] = 1;
        outs[63] = 62;
      end
      else begin
        valid[63] = 0;
        outs[63] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[63]) begin
      valid[64] = 1;
      outs[64] = outs[63];
    end
    else begin
      if (decode_signal[63]) begin
        valid[64] = 1;
        outs[64] = 63;
      end
      else begin
        valid[64] = 0;
        outs[64] = 0;
      end
    end
  end


endmodule // PriorityDecoder_0x2e5c0266b409153a

//-----------------------------------------------------------------------------
// CSRManager_0x68582ff11a9d1315
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.csr_manager {"interface": "op <C> (csr: Bits(12), rs1_is_x0: Bits(1), value: Bits(64), op: Bits(2)) -> (old: Bits(64), success: Bits(1))"}
// PyMTL: verilator_xinit = zeros
module CSRManager_0x68582ff11a9d1315
(
  input  logic [   0:0] clk,
  output logic  [   0:0] debug_recv_call,
  input  logic [  63:0] debug_recv_msg,
  input  logic [   0:0] debug_recv_rdy,
  output logic  [   0:0] debug_send_call,
  output logic  [  63:0] debug_send_msg,
  input  logic [   0:0] debug_send_rdy,
  input  logic [   0:0] op_call,
  input  logic [  11:0] op_csr,
  output logic  [  63:0] op_old,
  input  logic [   1:0] op_op,
  input  logic [   0:0] op_rs1_is_x0,
  output logic  [   0:0] op_success,
  input  logic [  63:0] op_value,
  input  logic [   0:0] reset
);

  // register declarations
  logic    [   0:0] temp_debug_recv_call;
  logic    [   0:0] temp_debug_send_call;
  logic    [  63:0] temp_debug_send_msg;
  logic    [  63:0] temp_op_old;
  logic    [   0:0] temp_op_success;

  // localparam declarations
  localparam CSR_FUNC_READ_WRITE = 2'd0;
  localparam mngr2proc = 12'd4032;
  localparam proc2mngr = 12'd1984;



  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_op():
  //       s.temp_debug_recv_call.v = 0
  //
  //       s.temp_debug_send_call.v = 0
  //       s.temp_debug_send_msg.v = 0
  //
  //       s.temp_op_success.v = 0
  //       s.temp_op_old.v = 0
  //
  //       if s.op_call:
  //         if s.op_csr == CsrRegisters.proc2mngr:
  //           if s.op_op == CsrFunc.CSR_FUNC_READ_WRITE and s.debug_send_rdy:
  //             s.temp_debug_send_call.v = 1
  //             s.temp_debug_send_msg.v = s.op_value
  //
  //             s.temp_op_success.v = 1
  //             s.temp_op_old.v = 0
  //         elif s.op_csr == CsrRegisters.mngr2proc:
  //           if s.op_op != CsrFunc.CSR_FUNC_READ_WRITE and s.debug_recv_rdy and s.op_rs1_is_x0:
  //             s.temp_debug_recv_call.v = 1
  //
  //             s.temp_op_success.v = 1
  //             s.temp_op_old.v = s.debug_recv_msg
  //
  //       s.debug_recv_call.v = s.temp_debug_recv_call
  //       s.debug_send_call.v = s.temp_debug_send_call
  //       s.debug_send_msg.v = s.temp_debug_send_msg
  //       s.op_success.v = s.temp_op_success
  //       s.op_old.v = s.temp_op_old

  // logic for handle_op()
  always @ (*) begin
    temp_debug_recv_call = 0;
    temp_debug_send_call = 0;
    temp_debug_send_msg = 0;
    temp_op_success = 0;
    temp_op_old = 0;
    if (op_call) begin
      if ((op_csr == proc2mngr)) begin
        if (((op_op == CSR_FUNC_READ_WRITE)&&debug_send_rdy)) begin
          temp_debug_send_call = 1;
          temp_debug_send_msg = op_value;
          temp_op_success = 1;
          temp_op_old = 0;
        end
        else begin
        end
      end
      else begin
        if ((op_csr == mngr2proc)) begin
          if (((op_op != CSR_FUNC_READ_WRITE)&&debug_recv_rdy&&op_rs1_is_x0)) begin
            temp_debug_recv_call = 1;
            temp_op_success = 1;
            temp_op_old = debug_recv_msg;
          end
          else begin
          end
        end
        else begin
        end
      end
    end
    else begin
    end
    debug_recv_call = temp_debug_recv_call;
    debug_send_call = temp_debug_send_call;
    debug_send_msg = temp_debug_send_msg;
    op_success = temp_op_success;
    op_old = temp_op_old;
  end


endmodule // CSRManager_0x68582ff11a9d1315

//-----------------------------------------------------------------------------
// GS14LWritebackStage23LWritebackDropController_0x4a102c6dab533550
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"args": ["process <C> (in_: Bits(146)) -> (accepted: Bits(1), out: Bits(142))"], "kwargs": {}}
// PyMTL: verilator_xinit = zeros
module GS14LWritebackStage23LWritebackDropController_0x4a102c6dab533550
(
  input  logic [   0:0] clk,
  output logic [   0:0] dataflow_write_call,
  output logic [   5:0] dataflow_write_tag,
  output logic [  63:0] dataflow_write_value,
  input  logic [ 145:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 141:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // pipeline_stage temporaries
  logic   [   0:0] pipeline_stage$check_keep;
  logic   [ 145:0] pipeline_stage$in_peek_msg;
  logic   [   0:0] pipeline_stage$clk;
  logic   [   4:0] pipeline_stage$kill_notify_msg;
  logic   [   0:0] pipeline_stage$in_peek_rdy;
  logic   [   0:0] pipeline_stage$process_accepted;
  logic   [ 141:0] pipeline_stage$check_out;
  logic   [   0:0] pipeline_stage$reset;
  logic   [ 141:0] pipeline_stage$process_out;
  logic   [   0:0] pipeline_stage$take_call;
  logic   [   0:0] pipeline_stage$process_call;
  logic   [ 141:0] pipeline_stage$check_in_;
  logic   [ 141:0] pipeline_stage$peek_msg;
  logic   [   4:0] pipeline_stage$check_msg;
  logic   [   0:0] pipeline_stage$in_take_call;
  logic   [   0:0] pipeline_stage$peek_rdy;
  logic   [ 145:0] pipeline_stage$process_in_;

  PipelineStage_0x6942ffa265da2f08 pipeline_stage
  (
    .check_keep       ( pipeline_stage$check_keep ),
    .in_peek_msg      ( pipeline_stage$in_peek_msg ),
    .clk              ( pipeline_stage$clk ),
    .kill_notify_msg  ( pipeline_stage$kill_notify_msg ),
    .in_peek_rdy      ( pipeline_stage$in_peek_rdy ),
    .process_accepted ( pipeline_stage$process_accepted ),
    .check_out        ( pipeline_stage$check_out ),
    .reset            ( pipeline_stage$reset ),
    .process_out      ( pipeline_stage$process_out ),
    .take_call        ( pipeline_stage$take_call ),
    .process_call     ( pipeline_stage$process_call ),
    .check_in_        ( pipeline_stage$check_in_ ),
    .peek_msg         ( pipeline_stage$peek_msg ),
    .check_msg        ( pipeline_stage$check_msg ),
    .in_take_call     ( pipeline_stage$in_take_call ),
    .peek_rdy         ( pipeline_stage$peek_rdy ),
    .process_in_      ( pipeline_stage$process_in_ )
  );

  // drop_controller temporaries
  logic   [   0:0] drop_controller$clk;
  logic   [ 141:0] drop_controller$check_in_;
  logic   [   4:0] drop_controller$check_msg;
  logic   [   0:0] drop_controller$reset;
  logic   [   0:0] drop_controller$check_keep;
  logic   [ 141:0] drop_controller$check_out;

  PipelineKillDropController_0x6535c882219b5c15 drop_controller
  (
    .clk        ( drop_controller$clk ),
    .check_in_  ( drop_controller$check_in_ ),
    .check_msg  ( drop_controller$check_msg ),
    .reset      ( drop_controller$reset ),
    .check_keep ( drop_controller$check_keep ),
    .check_out  ( drop_controller$check_out )
  );

  // stage temporaries
  logic   [   0:0] stage$process_call;
  logic   [   0:0] stage$clk;
  logic   [   0:0] stage$reset;
  logic   [ 145:0] stage$process_in_;
  logic   [   0:0] stage$dataflow_write_call;
  logic   [   0:0] stage$process_accepted;
  logic   [   5:0] stage$dataflow_write_tag;
  logic   [  63:0] stage$dataflow_write_value;
  logic   [ 141:0] stage$process_out;

  WritebackStage_0x620bfcc35a926f41 stage
  (
    .process_call         ( stage$process_call ),
    .clk                  ( stage$clk ),
    .reset                ( stage$reset ),
    .process_in_          ( stage$process_in_ ),
    .dataflow_write_call  ( stage$dataflow_write_call ),
    .process_accepted     ( stage$process_accepted ),
    .dataflow_write_tag   ( stage$dataflow_write_tag ),
    .dataflow_write_value ( stage$dataflow_write_value ),
    .process_out          ( stage$process_out )
  );

  // signal connections
  assign dataflow_write_call             = stage$dataflow_write_call;
  assign dataflow_write_tag              = stage$dataflow_write_tag;
  assign dataflow_write_value            = stage$dataflow_write_value;
  assign drop_controller$check_in_       = pipeline_stage$check_in_;
  assign drop_controller$check_msg       = pipeline_stage$check_msg;
  assign drop_controller$clk             = clk;
  assign drop_controller$reset           = reset;
  assign in_take_call                    = pipeline_stage$in_take_call;
  assign peek_msg                        = pipeline_stage$peek_msg;
  assign peek_rdy                        = pipeline_stage$peek_rdy;
  assign pipeline_stage$check_keep       = drop_controller$check_keep;
  assign pipeline_stage$check_out        = drop_controller$check_out;
  assign pipeline_stage$clk              = clk;
  assign pipeline_stage$in_peek_msg      = in_peek_msg;
  assign pipeline_stage$in_peek_rdy      = in_peek_rdy;
  assign pipeline_stage$kill_notify_msg  = kill_notify_msg;
  assign pipeline_stage$process_accepted = stage$process_accepted;
  assign pipeline_stage$process_out      = stage$process_out;
  assign pipeline_stage$reset            = reset;
  assign pipeline_stage$take_call        = take_call;
  assign stage$clk                       = clk;
  assign stage$process_call              = pipeline_stage$process_call;
  assign stage$process_in_               = pipeline_stage$process_in_;
  assign stage$reset                     = reset;



endmodule // GS14LWritebackStage23LWritebackDropController_0x4a102c6dab533550

//-----------------------------------------------------------------------------
// PipelineStage_0x6942ffa265da2f08
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.pipeline_stage {"In": 146, "Intermediate": null, "interface": "kill_notify (msg: Bits(5)) -> (); peek <R> () -> (msg: Bits(142)); take <C> () -> ()"}
// PyMTL: verilator_xinit = zeros
module PipelineStage_0x6942ffa265da2f08
(
  output logic [ 141:0] check_in_,
  input  logic [   0:0] check_keep,
  output logic [   4:0] check_msg,
  input  logic [ 141:0] check_out,
  input  logic [   0:0] clk,
  input  logic [ 145:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  output logic [ 141:0] peek_msg,
  output logic [   0:0] peek_rdy,
  input  logic [   0:0] process_accepted,
  output logic [   0:0] process_call,
  output logic [ 145:0] process_in_,
  input  logic [ 141:0] process_out,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // logic declarations
  logic   [   0:0] output_clear;
  logic   [   0:0] input_available;


  // register declarations
  logic    [   0:0] advance;
  logic    [   0:0] taking;

  // vvm temporaries
  logic   [   0:0] vvm$check_keep;
  logic   [   0:0] vvm$clk;
  logic   [   4:0] vvm$kill_notify_msg;
  logic   [ 141:0] vvm$add_msg;
  logic   [ 141:0] vvm$check_out;
  logic   [   0:0] vvm$reset;
  logic   [   0:0] vvm$add_call;
  logic   [   0:0] vvm$take_call;
  logic   [ 141:0] vvm$check_in_;
  logic   [ 141:0] vvm$peek_msg;
  logic   [   0:0] vvm$add_rdy;
  logic   [   4:0] vvm$check_msg;
  logic   [   0:0] vvm$peek_rdy;

  ValidValueManager_0xed9504a4389a8c9 vvm
  (
    .check_keep      ( vvm$check_keep ),
    .clk             ( vvm$clk ),
    .kill_notify_msg ( vvm$kill_notify_msg ),
    .add_msg         ( vvm$add_msg ),
    .check_out       ( vvm$check_out ),
    .reset           ( vvm$reset ),
    .add_call        ( vvm$add_call ),
    .take_call       ( vvm$take_call ),
    .check_in_       ( vvm$check_in_ ),
    .peek_msg        ( vvm$peek_msg ),
    .add_rdy         ( vvm$add_rdy ),
    .check_msg       ( vvm$check_msg ),
    .peek_rdy        ( vvm$peek_rdy )
  );

  // signal connections
  assign check_in_           = vvm$check_in_;
  assign check_msg           = vvm$check_msg;
  assign in_take_call        = taking;
  assign input_available     = in_peek_rdy;
  assign output_clear        = vvm$add_rdy;
  assign peek_msg            = vvm$peek_msg;
  assign peek_rdy            = vvm$peek_rdy;
  assign process_call        = advance;
  assign process_in_         = in_peek_msg;
  assign vvm$add_call        = taking;
  assign vvm$add_msg         = process_out;
  assign vvm$check_keep      = check_keep;
  assign vvm$check_out       = check_out;
  assign vvm$clk             = clk;
  assign vvm$kill_notify_msg = kill_notify_msg;
  assign vvm$reset           = reset;
  assign vvm$take_call       = take_call;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_taking():
  //       s.taking.v = s.advance & s.process_accepted

  // logic for handle_taking()
  always @ (*) begin
    taking = (advance&process_accepted);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_advance():
  //       s.advance.v = s.output_clear and s.input_available

  // logic for handle_advance()
  always @ (*) begin
    advance = (output_clear&&input_available);
  end


endmodule // PipelineStage_0x6942ffa265da2f08

//-----------------------------------------------------------------------------
// WritebackStage_0x620bfcc35a926f41
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.backend.writeback {"interface": "process <C> (in_: Bits(146)) -> (accepted: Bits(1), out: Bits(142))"}
// PyMTL: verilator_xinit = zeros
module WritebackStage_0x620bfcc35a926f41
(
  input  logic [   0:0] clk,
  output logic  [   0:0] dataflow_write_call,
  output logic  [   5:0] dataflow_write_tag,
  output logic  [  63:0] dataflow_write_value,
  output logic [   0:0] process_accepted,
  input  logic [   0:0] process_call,
  input  logic [ 145:0] process_in_,
  output logic  [ 141:0] process_out,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam PIPELINE_MSG_STATUS_VALID = 2'd0;

  // signal connections
  assign process_accepted = 1'd1;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute():
  //       s.process_out.v = 0
  //       s.process_out.hdr.v = s.process_in_.hdr
  //
  //       s.dataflow_write_call.v = 0
  //       s.dataflow_write_tag.v = 0
  //       s.dataflow_write_value.v = 0
  //
  //       if s.process_call:
  //         if s.process_in_.hdr_status == PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID:
  //           s.process_out.rd_val_pair.v = s.process_in_.rd_val_pair
  //
  //           # write the data if the destination is valid
  //           s.dataflow_write_call.v = s.process_in_.rd_val
  //           s.dataflow_write_tag.v = s.process_in_.rd
  //           s.dataflow_write_value.v = s.process_in_.result
  //         else:
  //           s.process_out.exception_info.v = s.process_in_.exception_info

  // logic for compute()
  always @ (*) begin
    process_out = 0;
    process_out[(74)-1:0] = process_in_[(74)-1:0];
    dataflow_write_call = 0;
    dataflow_write_tag = 0;
    dataflow_write_value = 0;
    if (process_call) begin
      if ((process_in_[(2)-1:0] == PIPELINE_MSG_STATUS_VALID)) begin
        process_out[(81)-1:74] = process_in_[(81)-1:74];
        dataflow_write_call = process_in_[(75)-1:74];
        dataflow_write_tag = process_in_[(81)-1:75];
        dataflow_write_value = process_in_[(146)-1:82];
      end
      else begin
        process_out[(142)-1:74] = process_in_[(142)-1:74];
      end
    end
    else begin
    end
  end


endmodule // WritebackStage_0x620bfcc35a926f41

//-----------------------------------------------------------------------------
// PipeSelector_0x7f9520fbc84f298e
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.backend.pipe_selector {}
// PyMTL: verilator_xinit = zeros
module PipeSelector_0x7f9520fbc84f298e
(
  output logic [ 250:0] alu_peek_msg,
  output logic [   0:0] alu_peek_rdy,
  input  logic [   0:0] alu_take_call,
  output logic [ 250:0] branch_peek_msg,
  output logic [   0:0] branch_peek_rdy,
  input  logic [   0:0] branch_take_call,
  input  logic [   0:0] clk,
  output logic [ 250:0] csr_peek_msg,
  output logic [   0:0] csr_peek_rdy,
  input  logic [   0:0] csr_take_call,
  input  logic [ 250:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   0:0] reset
);

  // splitter temporaries
  logic   [ 250:0] splitter$in_peek_msg;
  logic   [   0:0] splitter$branch_take_call;
  logic   [   0:0] splitter$alu_take_call;
  logic   [   0:0] splitter$clk;
  logic   [   0:0] splitter$in_peek_rdy;
  logic   [   1:0] splitter$sort_pipe;
  logic   [   0:0] splitter$reset;
  logic   [   0:0] splitter$csr_take_call;
  logic   [ 250:0] splitter$alu_peek_msg;
  logic   [   0:0] splitter$branch_peek_rdy;
  logic   [ 250:0] splitter$sort_msg;
  logic   [   0:0] splitter$alu_peek_rdy;
  logic   [ 250:0] splitter$branch_peek_msg;
  logic   [   0:0] splitter$in_take_call;
  logic   [   0:0] splitter$csr_peek_rdy;
  logic   [ 250:0] splitter$csr_peek_msg;

  PipelineSplitter_0x1033494f8d3884b8 splitter
  (
    .in_peek_msg      ( splitter$in_peek_msg ),
    .branch_take_call ( splitter$branch_take_call ),
    .alu_take_call    ( splitter$alu_take_call ),
    .clk              ( splitter$clk ),
    .in_peek_rdy      ( splitter$in_peek_rdy ),
    .sort_pipe        ( splitter$sort_pipe ),
    .reset            ( splitter$reset ),
    .csr_take_call    ( splitter$csr_take_call ),
    .alu_peek_msg     ( splitter$alu_peek_msg ),
    .branch_peek_rdy  ( splitter$branch_peek_rdy ),
    .sort_msg         ( splitter$sort_msg ),
    .alu_peek_rdy     ( splitter$alu_peek_rdy ),
    .branch_peek_msg  ( splitter$branch_peek_msg ),
    .in_take_call     ( splitter$in_take_call ),
    .csr_peek_rdy     ( splitter$csr_peek_rdy ),
    .csr_peek_msg     ( splitter$csr_peek_msg )
  );

  // controller temporaries
  logic   [   0:0] controller$clk;
  logic   [ 250:0] controller$sort_msg;
  logic   [   0:0] controller$reset;
  logic   [   1:0] controller$sort_pipe;

  PipeSelectorController_0x7f9520fbc84f298e controller
  (
    .clk       ( controller$clk ),
    .sort_msg  ( controller$sort_msg ),
    .reset     ( controller$reset ),
    .sort_pipe ( controller$sort_pipe )
  );

  // signal connections
  assign alu_peek_msg              = splitter$alu_peek_msg;
  assign alu_peek_rdy              = splitter$alu_peek_rdy;
  assign branch_peek_msg           = splitter$branch_peek_msg;
  assign branch_peek_rdy           = splitter$branch_peek_rdy;
  assign controller$clk            = clk;
  assign controller$reset          = reset;
  assign controller$sort_msg       = splitter$sort_msg;
  assign csr_peek_msg              = splitter$csr_peek_msg;
  assign csr_peek_rdy              = splitter$csr_peek_rdy;
  assign in_take_call              = splitter$in_take_call;
  assign splitter$alu_take_call    = alu_take_call;
  assign splitter$branch_take_call = branch_take_call;
  assign splitter$clk              = clk;
  assign splitter$csr_take_call    = csr_take_call;
  assign splitter$in_peek_msg      = in_peek_msg;
  assign splitter$in_peek_rdy      = in_peek_rdy;
  assign splitter$reset            = reset;
  assign splitter$sort_pipe        = controller$sort_pipe;



endmodule // PipeSelector_0x7f9520fbc84f298e

//-----------------------------------------------------------------------------
// PipelineSplitter_0x1033494f8d3884b8
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.pipeline_splitter {"interface": "csr_peek <R> () -> (msg: Bits(251)); csr_take <C> () -> (); alu_peek <R> () -> (msg: Bits(251)); alu_take <C> () -> (); branch_peek <R> () -> (msg: Bits(251)); branch_take <C> () -> ()"}
// PyMTL: verilator_xinit = zeros
module PipelineSplitter_0x1033494f8d3884b8
(
  output logic [ 250:0] alu_peek_msg,
  output logic [   0:0] alu_peek_rdy,
  input  logic [   0:0] alu_take_call,
  output logic [ 250:0] branch_peek_msg,
  output logic [   0:0] branch_peek_rdy,
  input  logic [   0:0] branch_take_call,
  input  logic [   0:0] clk,
  output logic [ 250:0] csr_peek_msg,
  output logic [   0:0] csr_peek_rdy,
  input  logic [   0:0] csr_take_call,
  input  logic [ 250:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   0:0] reset,
  output logic [ 250:0] sort_msg,
  input  logic [   1:0] sort_pipe
);

  // logic declarations
  logic   [   0:0] effective_call;
  logic   [   0:0] rdy_array$000;
  logic   [   0:0] rdy_array$001;
  logic   [   0:0] rdy_array$002;


  // take_mux temporaries
  logic   [   0:0] take_mux$mux_in_$000;
  logic   [   0:0] take_mux$mux_in_$001;
  logic   [   0:0] take_mux$mux_in_$002;
  logic   [   0:0] take_mux$clk;
  logic   [   0:0] take_mux$reset;
  logic   [   1:0] take_mux$mux_select;
  logic   [   0:0] take_mux$mux_out;

  Mux_0x183cf582fc9c6432 take_mux
  (
    .mux_in_$000 ( take_mux$mux_in_$000 ),
    .mux_in_$001 ( take_mux$mux_in_$001 ),
    .mux_in_$002 ( take_mux$mux_in_$002 ),
    .clk         ( take_mux$clk ),
    .reset       ( take_mux$reset ),
    .mux_select  ( take_mux$mux_select ),
    .mux_out     ( take_mux$mux_out )
  );

  // signal connections
  assign alu_peek_msg         = in_peek_msg;
  assign alu_peek_rdy         = rdy_array$001;
  assign branch_peek_msg      = in_peek_msg;
  assign branch_peek_rdy      = rdy_array$002;
  assign csr_peek_msg         = in_peek_msg;
  assign csr_peek_rdy         = rdy_array$000;
  assign in_take_call         = take_mux$mux_out;
  assign sort_msg             = in_peek_msg;
  assign take_mux$clk         = clk;
  assign take_mux$mux_in_$000 = csr_take_call;
  assign take_mux$mux_in_$001 = alu_take_call;
  assign take_mux$mux_in_$002 = branch_take_call;
  assign take_mux$mux_select  = sort_pipe;
  assign take_mux$reset       = reset;

  // array declarations
  logic    [   0:0] rdy_array[0:2];
  assign rdy_array$000 = rdy_array[  0];
  assign rdy_array$001 = rdy_array[  1];
  assign rdy_array$002 = rdy_array[  2];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_rdy(i=i):
  //         s.rdy_array[i].v = (s.sort_pipe == i) and s.in_peek_rdy

  // logic for handle_rdy()
  always @ (*) begin
    rdy_array[0] = ((sort_pipe == 0)&&in_peek_rdy);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_rdy(i=i):
  //         s.rdy_array[i].v = (s.sort_pipe == i) and s.in_peek_rdy

  // logic for handle_rdy()
  always @ (*) begin
    rdy_array[1] = ((sort_pipe == 1)&&in_peek_rdy);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_rdy(i=i):
  //         s.rdy_array[i].v = (s.sort_pipe == i) and s.in_peek_rdy

  // logic for handle_rdy()
  always @ (*) begin
    rdy_array[2] = ((sort_pipe == 2)&&in_peek_rdy);
  end


endmodule // PipelineSplitter_0x1033494f8d3884b8

//-----------------------------------------------------------------------------
// Mux_0x183cf582fc9c6432
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.mux {"dtype": 1, "nports": 3}
// PyMTL: verilator_xinit = zeros
module Mux_0x183cf582fc9c6432
(
  input  logic [   0:0] clk,
  input  logic [   0:0] mux_in_$000,
  input  logic [   0:0] mux_in_$001,
  input  logic [   0:0] mux_in_$002,
  output logic  [   0:0] mux_out,
  input  logic [   1:0] mux_select,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nports = 3;


  // array declarations
  logic   [   0:0] mux_in_[0:2];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def select():
  //       assert s.mux_select < nports
  //       s.mux_out.v = s.mux_in_[s.mux_select]

  // logic for select()
  always @ (*) begin
    mux_out = mux_in_[mux_select];
  end


endmodule // Mux_0x183cf582fc9c6432

//-----------------------------------------------------------------------------
// PipeSelectorController_0x7f9520fbc84f298e
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.backend.pipe_selector {}
// PyMTL: verilator_xinit = zeros
module PipeSelectorController_0x7f9520fbc84f298e
(
  input  logic [   0:0] clk,
  input  logic [   0:0] reset,
  input  logic [ 250:0] sort_msg,
  output logic  [   1:0] sort_pipe
);

  // localparam declarations
  localparam OP_CLASS_ALU = 3'd0;
  localparam OP_CLASS_BRANCH = 3'd2;
  localparam OP_CLASS_CSR = 3'd3;
  localparam PIPELINE_MSG_STATUS_VALID = 2'd0;



  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_sort():
  //       if s.sort_msg.hdr_status != PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID:
  //         s.sort_pipe.v = 0  # CSR pipe
  //       elif s.sort_msg.op_class == OpClass.OP_CLASS_CSR:
  //         s.sort_pipe.v = 0  # CSR pipe
  //       elif s.sort_msg.op_class == OpClass.OP_CLASS_ALU:
  //         s.sort_pipe.v = 1  # ALU pipe
  //       elif s.sort_msg.op_class == OpClass.OP_CLASS_BRANCH:
  //         s.sort_pipe.v = 2  # Branch pipe
  //       else:
  //         s.sort_pipe.v = 0  # Error CSR pipe

  // logic for handle_sort()
  always @ (*) begin
    if ((sort_msg[(2)-1:0] != PIPELINE_MSG_STATUS_VALID)) begin
      sort_pipe = 0;
    end
    else begin
      if ((sort_msg[(236)-1:233] == OP_CLASS_CSR)) begin
        sort_pipe = 0;
      end
      else begin
        if ((sort_msg[(236)-1:233] == OP_CLASS_ALU)) begin
          sort_pipe = 1;
        end
        else begin
          if ((sort_msg[(236)-1:233] == OP_CLASS_BRANCH)) begin
            sort_pipe = 2;
          end
          else begin
            sort_pipe = 0;
          end
        end
      end
    end
  end


endmodule // PipeSelectorController_0x7f9520fbc84f298e

//-----------------------------------------------------------------------------
// DataFlowManager_0x54912d9190dab9c9
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.dataflow {"dflow_interface": "is_ready[2] (tag: Bits(6)) -> (ready: Bits(1)); write[1] <C> (tag: Bits(6), value: Bits(64)) -> (); get_updated () -> (mask: Bits(64)); get_src[2] (areg: Bits(5)) -> (preg: Bits(6)); get_dst[1] <CR> (areg: Bits(5)) -> (preg: Bits(6)); commit[1] <C> (tag: Bits(6)) -> (); read[2] (tag: Bits(6)) -> (value: Bits(64)); snapshot <CR> () -> (id_: Bits(1)); free_snapshot <C> (id_: Bits(1)) -> (); restore <C> (source_id: Bits(1)) -> (); rollback <C> () -> ()"}
// PyMTL: verilator_xinit = zeros
module DataFlowManager_0x54912d9190dab9c9
(
  input  logic [   0:0] clk,
  input  logic [   0:0] commit_call$000,
  input  logic [   5:0] commit_tag$000,
  input  logic [   0:0] free_snapshot_call,
  input  logic [   0:0] free_snapshot_id_,
  input  logic [   4:0] get_dst_areg$000,
  input  logic [   0:0] get_dst_call$000,
  output logic [   5:0] get_dst_preg$000,
  output logic [   0:0] get_dst_rdy$000,
  input  logic [   4:0] get_src_areg$000,
  input  logic [   4:0] get_src_areg$001,
  output logic [   5:0] get_src_preg$000,
  output logic [   5:0] get_src_preg$001,
  output logic [  63:0] get_updated_mask,
  output logic [   0:0] is_ready_ready$000,
  output logic [   0:0] is_ready_ready$001,
  input  logic [   5:0] is_ready_tag$000,
  input  logic [   5:0] is_ready_tag$001,
  input  logic [   5:0] read_tag$000,
  input  logic [   5:0] read_tag$001,
  output logic [  63:0] read_value$000,
  output logic [  63:0] read_value$001,
  input  logic [   0:0] reset,
  input  logic [   0:0] restore_call,
  input  logic [   0:0] restore_source_id,
  input  logic [   0:0] rollback_call,
  input  logic [   0:0] snapshot_call,
  output logic [   0:0] snapshot_id_,
  output logic [   0:0] snapshot_rdy,
  input  logic [   0:0] write_call$000,
  input  logic [   5:0] write_tag$000,
  input  logic [  63:0] write_value$000
);

  // logic declarations
  logic   [  63:0] get_updated_incremental_masks$000;
  logic   [  63:0] get_updated_incremental_masks$001;
  logic   [   0:0] is_ready_is_zero_tag$000;
  logic   [   0:0] is_ready_is_zero_tag$001;
  logic   [   0:0] read_is_zero_tag$000;
  logic   [   0:0] read_is_zero_tag$001;
  logic   [   0:0] is_write_not_zero_tag$000;
  logic   [   0:0] is_commit_not_zero_tag$000;
  logic   [   0:0] get_dst_need_writeback$000;


  // register declarations
  logic    [  62:0] free_regs$set_state;

  // localparam declarations
  localparam ZERO_TAG = 6'd63;

  // snapshot_allocator temporaries
  logic   [   1:0] snapshot_allocator$set_state;
  logic   [   0:0] snapshot_allocator$revert_allocs_call;
  logic   [   0:0] snapshot_allocator$set_call;
  logic   [   0:0] snapshot_allocator$revert_allocs_source_id;
  logic   [   0:0] snapshot_allocator$clk;
  logic   [   0:0] snapshot_allocator$free_call$000;
  logic   [   0:0] snapshot_allocator$reset_alloc_tracking_call;
  logic   [   0:0] snapshot_allocator$reset_alloc_tracking_target_id;
  logic   [   0:0] snapshot_allocator$alloc_call$000;
  logic   [   0:0] snapshot_allocator$reset;
  logic   [   0:0] snapshot_allocator$free_index$000;
  logic   [   1:0] snapshot_allocator$alloc_mask$000;
  logic   [   0:0] snapshot_allocator$alloc_rdy$000;
  logic   [   0:0] snapshot_allocator$alloc_index$000;

  SnapshottingFreeList_0x64ee202bb6767a5b snapshot_allocator
  (
    .set_state                      ( snapshot_allocator$set_state ),
    .revert_allocs_call             ( snapshot_allocator$revert_allocs_call ),
    .set_call                       ( snapshot_allocator$set_call ),
    .revert_allocs_source_id        ( snapshot_allocator$revert_allocs_source_id ),
    .clk                            ( snapshot_allocator$clk ),
    .free_call$000                  ( snapshot_allocator$free_call$000 ),
    .reset_alloc_tracking_call      ( snapshot_allocator$reset_alloc_tracking_call ),
    .reset_alloc_tracking_target_id ( snapshot_allocator$reset_alloc_tracking_target_id ),
    .alloc_call$000                 ( snapshot_allocator$alloc_call$000 ),
    .reset                          ( snapshot_allocator$reset ),
    .free_index$000                 ( snapshot_allocator$free_index$000 ),
    .alloc_mask$000                 ( snapshot_allocator$alloc_mask$000 ),
    .alloc_rdy$000                  ( snapshot_allocator$alloc_rdy$000 ),
    .alloc_index$000                ( snapshot_allocator$alloc_index$000 )
  );

  // ready_table temporaries
  logic   [   0:0] ready_table$clk;
  logic   [   5:0] ready_table$write_addr$000;
  logic   [   5:0] ready_table$write_addr$001;
  logic   [   5:0] ready_table$read_addr$000;
  logic   [   5:0] ready_table$read_addr$001;
  logic   [   0:0] ready_table$write_call$000;
  logic   [   0:0] ready_table$write_call$001;
  logic   [   0:0] ready_table$write_data$000;
  logic   [   0:0] ready_table$write_data$001;
  logic   [   0:0] ready_table$reset;
  logic   [   0:0] ready_table$read_data$000;
  logic   [   0:0] ready_table$read_data$001;

  AsynchronousRAM_0x49021b1555bbbcb6 ready_table
  (
    .clk            ( ready_table$clk ),
    .write_addr$000 ( ready_table$write_addr$000 ),
    .write_addr$001 ( ready_table$write_addr$001 ),
    .read_addr$000  ( ready_table$read_addr$000 ),
    .read_addr$001  ( ready_table$read_addr$001 ),
    .write_call$000 ( ready_table$write_call$000 ),
    .write_call$001 ( ready_table$write_call$001 ),
    .write_data$000 ( ready_table$write_data$000 ),
    .write_data$001 ( ready_table$write_data$001 ),
    .reset          ( ready_table$reset ),
    .read_data$000  ( ready_table$read_data$000 ),
    .read_data$001  ( ready_table$read_data$001 )
  );

  // read_muxes_ready$000 temporaries
  logic   [   0:0] read_muxes_ready$000$mux_in_$000;
  logic   [   0:0] read_muxes_ready$000$mux_in_$001;
  logic   [   0:0] read_muxes_ready$000$clk;
  logic   [   0:0] read_muxes_ready$000$reset;
  logic   [   0:0] read_muxes_ready$000$mux_select;
  logic   [   0:0] read_muxes_ready$000$mux_out;

  Mux_0x183cf582fc8d227d read_muxes_ready$000
  (
    .mux_in_$000 ( read_muxes_ready$000$mux_in_$000 ),
    .mux_in_$001 ( read_muxes_ready$000$mux_in_$001 ),
    .clk         ( read_muxes_ready$000$clk ),
    .reset       ( read_muxes_ready$000$reset ),
    .mux_select  ( read_muxes_ready$000$mux_select ),
    .mux_out     ( read_muxes_ready$000$mux_out )
  );

  // read_muxes_ready$001 temporaries
  logic   [   0:0] read_muxes_ready$001$mux_in_$000;
  logic   [   0:0] read_muxes_ready$001$mux_in_$001;
  logic   [   0:0] read_muxes_ready$001$clk;
  logic   [   0:0] read_muxes_ready$001$reset;
  logic   [   0:0] read_muxes_ready$001$mux_select;
  logic   [   0:0] read_muxes_ready$001$mux_out;

  Mux_0x183cf582fc8d227d read_muxes_ready$001
  (
    .mux_in_$000 ( read_muxes_ready$001$mux_in_$000 ),
    .mux_in_$001 ( read_muxes_ready$001$mux_in_$001 ),
    .clk         ( read_muxes_ready$001$clk ),
    .reset       ( read_muxes_ready$001$reset ),
    .mux_select  ( read_muxes_ready$001$mux_select ),
    .mux_out     ( read_muxes_ready$001$mux_out )
  );

  // arch_used_pregs_packer temporaries
  logic   [   0:0] arch_used_pregs_packer$clk;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$000;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$001;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$002;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$003;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$004;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$005;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$006;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$007;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$008;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$009;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$010;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$011;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$012;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$013;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$014;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$015;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$016;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$017;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$018;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$019;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$020;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$021;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$022;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$023;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$024;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$025;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$026;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$027;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$028;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$029;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$030;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$031;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$032;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$033;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$034;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$035;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$036;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$037;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$038;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$039;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$040;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$041;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$042;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$043;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$044;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$045;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$046;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$047;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$048;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$049;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$050;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$051;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$052;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$053;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$054;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$055;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$056;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$057;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$058;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$059;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$060;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$061;
  logic   [   0:0] arch_used_pregs_packer$pack_in_$062;
  logic   [   0:0] arch_used_pregs_packer$reset;
  logic   [  62:0] arch_used_pregs_packer$pack_packed;

  Packer_0x5417ceb8bd59f204 arch_used_pregs_packer
  (
    .clk          ( arch_used_pregs_packer$clk ),
    .pack_in_$000 ( arch_used_pregs_packer$pack_in_$000 ),
    .pack_in_$001 ( arch_used_pregs_packer$pack_in_$001 ),
    .pack_in_$002 ( arch_used_pregs_packer$pack_in_$002 ),
    .pack_in_$003 ( arch_used_pregs_packer$pack_in_$003 ),
    .pack_in_$004 ( arch_used_pregs_packer$pack_in_$004 ),
    .pack_in_$005 ( arch_used_pregs_packer$pack_in_$005 ),
    .pack_in_$006 ( arch_used_pregs_packer$pack_in_$006 ),
    .pack_in_$007 ( arch_used_pregs_packer$pack_in_$007 ),
    .pack_in_$008 ( arch_used_pregs_packer$pack_in_$008 ),
    .pack_in_$009 ( arch_used_pregs_packer$pack_in_$009 ),
    .pack_in_$010 ( arch_used_pregs_packer$pack_in_$010 ),
    .pack_in_$011 ( arch_used_pregs_packer$pack_in_$011 ),
    .pack_in_$012 ( arch_used_pregs_packer$pack_in_$012 ),
    .pack_in_$013 ( arch_used_pregs_packer$pack_in_$013 ),
    .pack_in_$014 ( arch_used_pregs_packer$pack_in_$014 ),
    .pack_in_$015 ( arch_used_pregs_packer$pack_in_$015 ),
    .pack_in_$016 ( arch_used_pregs_packer$pack_in_$016 ),
    .pack_in_$017 ( arch_used_pregs_packer$pack_in_$017 ),
    .pack_in_$018 ( arch_used_pregs_packer$pack_in_$018 ),
    .pack_in_$019 ( arch_used_pregs_packer$pack_in_$019 ),
    .pack_in_$020 ( arch_used_pregs_packer$pack_in_$020 ),
    .pack_in_$021 ( arch_used_pregs_packer$pack_in_$021 ),
    .pack_in_$022 ( arch_used_pregs_packer$pack_in_$022 ),
    .pack_in_$023 ( arch_used_pregs_packer$pack_in_$023 ),
    .pack_in_$024 ( arch_used_pregs_packer$pack_in_$024 ),
    .pack_in_$025 ( arch_used_pregs_packer$pack_in_$025 ),
    .pack_in_$026 ( arch_used_pregs_packer$pack_in_$026 ),
    .pack_in_$027 ( arch_used_pregs_packer$pack_in_$027 ),
    .pack_in_$028 ( arch_used_pregs_packer$pack_in_$028 ),
    .pack_in_$029 ( arch_used_pregs_packer$pack_in_$029 ),
    .pack_in_$030 ( arch_used_pregs_packer$pack_in_$030 ),
    .pack_in_$031 ( arch_used_pregs_packer$pack_in_$031 ),
    .pack_in_$032 ( arch_used_pregs_packer$pack_in_$032 ),
    .pack_in_$033 ( arch_used_pregs_packer$pack_in_$033 ),
    .pack_in_$034 ( arch_used_pregs_packer$pack_in_$034 ),
    .pack_in_$035 ( arch_used_pregs_packer$pack_in_$035 ),
    .pack_in_$036 ( arch_used_pregs_packer$pack_in_$036 ),
    .pack_in_$037 ( arch_used_pregs_packer$pack_in_$037 ),
    .pack_in_$038 ( arch_used_pregs_packer$pack_in_$038 ),
    .pack_in_$039 ( arch_used_pregs_packer$pack_in_$039 ),
    .pack_in_$040 ( arch_used_pregs_packer$pack_in_$040 ),
    .pack_in_$041 ( arch_used_pregs_packer$pack_in_$041 ),
    .pack_in_$042 ( arch_used_pregs_packer$pack_in_$042 ),
    .pack_in_$043 ( arch_used_pregs_packer$pack_in_$043 ),
    .pack_in_$044 ( arch_used_pregs_packer$pack_in_$044 ),
    .pack_in_$045 ( arch_used_pregs_packer$pack_in_$045 ),
    .pack_in_$046 ( arch_used_pregs_packer$pack_in_$046 ),
    .pack_in_$047 ( arch_used_pregs_packer$pack_in_$047 ),
    .pack_in_$048 ( arch_used_pregs_packer$pack_in_$048 ),
    .pack_in_$049 ( arch_used_pregs_packer$pack_in_$049 ),
    .pack_in_$050 ( arch_used_pregs_packer$pack_in_$050 ),
    .pack_in_$051 ( arch_used_pregs_packer$pack_in_$051 ),
    .pack_in_$052 ( arch_used_pregs_packer$pack_in_$052 ),
    .pack_in_$053 ( arch_used_pregs_packer$pack_in_$053 ),
    .pack_in_$054 ( arch_used_pregs_packer$pack_in_$054 ),
    .pack_in_$055 ( arch_used_pregs_packer$pack_in_$055 ),
    .pack_in_$056 ( arch_used_pregs_packer$pack_in_$056 ),
    .pack_in_$057 ( arch_used_pregs_packer$pack_in_$057 ),
    .pack_in_$058 ( arch_used_pregs_packer$pack_in_$058 ),
    .pack_in_$059 ( arch_used_pregs_packer$pack_in_$059 ),
    .pack_in_$060 ( arch_used_pregs_packer$pack_in_$060 ),
    .pack_in_$061 ( arch_used_pregs_packer$pack_in_$061 ),
    .pack_in_$062 ( arch_used_pregs_packer$pack_in_$062 ),
    .reset        ( arch_used_pregs_packer$reset ),
    .pack_packed  ( arch_used_pregs_packer$pack_packed )
  );

  // rename_table temporaries
  logic   [   0:0] rename_table$snapshot_call;
  logic   [   5:0] rename_table$set_in_$000;
  logic   [   5:0] rename_table$set_in_$001;
  logic   [   5:0] rename_table$set_in_$002;
  logic   [   5:0] rename_table$set_in_$003;
  logic   [   5:0] rename_table$set_in_$004;
  logic   [   5:0] rename_table$set_in_$005;
  logic   [   5:0] rename_table$set_in_$006;
  logic   [   5:0] rename_table$set_in_$007;
  logic   [   5:0] rename_table$set_in_$008;
  logic   [   5:0] rename_table$set_in_$009;
  logic   [   5:0] rename_table$set_in_$010;
  logic   [   5:0] rename_table$set_in_$011;
  logic   [   5:0] rename_table$set_in_$012;
  logic   [   5:0] rename_table$set_in_$013;
  logic   [   5:0] rename_table$set_in_$014;
  logic   [   5:0] rename_table$set_in_$015;
  logic   [   5:0] rename_table$set_in_$016;
  logic   [   5:0] rename_table$set_in_$017;
  logic   [   5:0] rename_table$set_in_$018;
  logic   [   5:0] rename_table$set_in_$019;
  logic   [   5:0] rename_table$set_in_$020;
  logic   [   5:0] rename_table$set_in_$021;
  logic   [   5:0] rename_table$set_in_$022;
  logic   [   5:0] rename_table$set_in_$023;
  logic   [   5:0] rename_table$set_in_$024;
  logic   [   5:0] rename_table$set_in_$025;
  logic   [   5:0] rename_table$set_in_$026;
  logic   [   5:0] rename_table$set_in_$027;
  logic   [   5:0] rename_table$set_in_$028;
  logic   [   5:0] rename_table$set_in_$029;
  logic   [   5:0] rename_table$set_in_$030;
  logic   [   5:0] rename_table$set_in_$031;
  logic   [   0:0] rename_table$update_call$000;
  logic   [   0:0] rename_table$set_call;
  logic   [   0:0] rename_table$restore_source_id;
  logic   [   0:0] rename_table$restore_call;
  logic   [   0:0] rename_table$clk;
  logic   [   4:0] rename_table$lookup_areg$000;
  logic   [   4:0] rename_table$lookup_areg$001;
  logic   [   4:0] rename_table$update_areg$000;
  logic   [   0:0] rename_table$snapshot_target_id;
  logic   [   5:0] rename_table$update_preg$000;
  logic   [   0:0] rename_table$reset;
  logic   [   5:0] rename_table$lookup_preg$000;
  logic   [   5:0] rename_table$lookup_preg$001;

  RenameTable_0x2b84c99320ad3cb1 rename_table
  (
    .snapshot_call      ( rename_table$snapshot_call ),
    .set_in_$000        ( rename_table$set_in_$000 ),
    .set_in_$001        ( rename_table$set_in_$001 ),
    .set_in_$002        ( rename_table$set_in_$002 ),
    .set_in_$003        ( rename_table$set_in_$003 ),
    .set_in_$004        ( rename_table$set_in_$004 ),
    .set_in_$005        ( rename_table$set_in_$005 ),
    .set_in_$006        ( rename_table$set_in_$006 ),
    .set_in_$007        ( rename_table$set_in_$007 ),
    .set_in_$008        ( rename_table$set_in_$008 ),
    .set_in_$009        ( rename_table$set_in_$009 ),
    .set_in_$010        ( rename_table$set_in_$010 ),
    .set_in_$011        ( rename_table$set_in_$011 ),
    .set_in_$012        ( rename_table$set_in_$012 ),
    .set_in_$013        ( rename_table$set_in_$013 ),
    .set_in_$014        ( rename_table$set_in_$014 ),
    .set_in_$015        ( rename_table$set_in_$015 ),
    .set_in_$016        ( rename_table$set_in_$016 ),
    .set_in_$017        ( rename_table$set_in_$017 ),
    .set_in_$018        ( rename_table$set_in_$018 ),
    .set_in_$019        ( rename_table$set_in_$019 ),
    .set_in_$020        ( rename_table$set_in_$020 ),
    .set_in_$021        ( rename_table$set_in_$021 ),
    .set_in_$022        ( rename_table$set_in_$022 ),
    .set_in_$023        ( rename_table$set_in_$023 ),
    .set_in_$024        ( rename_table$set_in_$024 ),
    .set_in_$025        ( rename_table$set_in_$025 ),
    .set_in_$026        ( rename_table$set_in_$026 ),
    .set_in_$027        ( rename_table$set_in_$027 ),
    .set_in_$028        ( rename_table$set_in_$028 ),
    .set_in_$029        ( rename_table$set_in_$029 ),
    .set_in_$030        ( rename_table$set_in_$030 ),
    .set_in_$031        ( rename_table$set_in_$031 ),
    .update_call$000    ( rename_table$update_call$000 ),
    .set_call           ( rename_table$set_call ),
    .restore_source_id  ( rename_table$restore_source_id ),
    .restore_call       ( rename_table$restore_call ),
    .clk                ( rename_table$clk ),
    .lookup_areg$000    ( rename_table$lookup_areg$000 ),
    .lookup_areg$001    ( rename_table$lookup_areg$001 ),
    .update_areg$000    ( rename_table$update_areg$000 ),
    .snapshot_target_id ( rename_table$snapshot_target_id ),
    .update_preg$000    ( rename_table$update_preg$000 ),
    .reset              ( rename_table$reset ),
    .lookup_preg$000    ( rename_table$lookup_preg$000 ),
    .lookup_preg$001    ( rename_table$lookup_preg$001 )
  );

  // inverse temporaries
  logic   [   0:0] inverse$clk;
  logic   [   5:0] inverse$write_addr$000;
  logic   [   5:0] inverse$read_addr$000;
  logic   [   0:0] inverse$write_call$000;
  logic   [   4:0] inverse$write_data$000;
  logic   [   0:0] inverse$reset;
  logic   [   4:0] inverse$read_data$000;

  AsynchronousRAM_0x6ff7d20a35694d13 inverse
  (
    .clk            ( inverse$clk ),
    .write_addr$000 ( inverse$write_addr$000 ),
    .read_addr$000  ( inverse$read_addr$000 ),
    .write_call$000 ( inverse$write_call$000 ),
    .write_data$000 ( inverse$write_data$000 ),
    .reset          ( inverse$reset ),
    .read_data$000  ( inverse$read_data$000 )
  );

  // areg_file temporaries
  logic   [   5:0] areg_file$set_in_$000;
  logic   [   5:0] areg_file$set_in_$001;
  logic   [   5:0] areg_file$set_in_$002;
  logic   [   5:0] areg_file$set_in_$003;
  logic   [   5:0] areg_file$set_in_$004;
  logic   [   5:0] areg_file$set_in_$005;
  logic   [   5:0] areg_file$set_in_$006;
  logic   [   5:0] areg_file$set_in_$007;
  logic   [   5:0] areg_file$set_in_$008;
  logic   [   5:0] areg_file$set_in_$009;
  logic   [   5:0] areg_file$set_in_$010;
  logic   [   5:0] areg_file$set_in_$011;
  logic   [   5:0] areg_file$set_in_$012;
  logic   [   5:0] areg_file$set_in_$013;
  logic   [   5:0] areg_file$set_in_$014;
  logic   [   5:0] areg_file$set_in_$015;
  logic   [   5:0] areg_file$set_in_$016;
  logic   [   5:0] areg_file$set_in_$017;
  logic   [   5:0] areg_file$set_in_$018;
  logic   [   5:0] areg_file$set_in_$019;
  logic   [   5:0] areg_file$set_in_$020;
  logic   [   5:0] areg_file$set_in_$021;
  logic   [   5:0] areg_file$set_in_$022;
  logic   [   5:0] areg_file$set_in_$023;
  logic   [   5:0] areg_file$set_in_$024;
  logic   [   5:0] areg_file$set_in_$025;
  logic   [   5:0] areg_file$set_in_$026;
  logic   [   5:0] areg_file$set_in_$027;
  logic   [   5:0] areg_file$set_in_$028;
  logic   [   5:0] areg_file$set_in_$029;
  logic   [   5:0] areg_file$set_in_$030;
  logic   [   5:0] areg_file$set_in_$031;
  logic   [   0:0] areg_file$set_call;
  logic   [   0:0] areg_file$clk;
  logic   [   4:0] areg_file$write_addr$000;
  logic   [   4:0] areg_file$read_addr$000;
  logic   [   0:0] areg_file$write_call$000;
  logic   [   5:0] areg_file$write_data$000;
  logic   [   0:0] areg_file$reset;
  logic   [   5:0] areg_file$read_data$000;
  logic   [   5:0] areg_file$dump_out$000;
  logic   [   5:0] areg_file$dump_out$001;
  logic   [   5:0] areg_file$dump_out$002;
  logic   [   5:0] areg_file$dump_out$003;
  logic   [   5:0] areg_file$dump_out$004;
  logic   [   5:0] areg_file$dump_out$005;
  logic   [   5:0] areg_file$dump_out$006;
  logic   [   5:0] areg_file$dump_out$007;
  logic   [   5:0] areg_file$dump_out$008;
  logic   [   5:0] areg_file$dump_out$009;
  logic   [   5:0] areg_file$dump_out$010;
  logic   [   5:0] areg_file$dump_out$011;
  logic   [   5:0] areg_file$dump_out$012;
  logic   [   5:0] areg_file$dump_out$013;
  logic   [   5:0] areg_file$dump_out$014;
  logic   [   5:0] areg_file$dump_out$015;
  logic   [   5:0] areg_file$dump_out$016;
  logic   [   5:0] areg_file$dump_out$017;
  logic   [   5:0] areg_file$dump_out$018;
  logic   [   5:0] areg_file$dump_out$019;
  logic   [   5:0] areg_file$dump_out$020;
  logic   [   5:0] areg_file$dump_out$021;
  logic   [   5:0] areg_file$dump_out$022;
  logic   [   5:0] areg_file$dump_out$023;
  logic   [   5:0] areg_file$dump_out$024;
  logic   [   5:0] areg_file$dump_out$025;
  logic   [   5:0] areg_file$dump_out$026;
  logic   [   5:0] areg_file$dump_out$027;
  logic   [   5:0] areg_file$dump_out$028;
  logic   [   5:0] areg_file$dump_out$029;
  logic   [   5:0] areg_file$dump_out$030;
  logic   [   5:0] areg_file$dump_out$031;

  RegisterFile_0x6ba986f42995f7d7 areg_file
  (
    .set_in_$000    ( areg_file$set_in_$000 ),
    .set_in_$001    ( areg_file$set_in_$001 ),
    .set_in_$002    ( areg_file$set_in_$002 ),
    .set_in_$003    ( areg_file$set_in_$003 ),
    .set_in_$004    ( areg_file$set_in_$004 ),
    .set_in_$005    ( areg_file$set_in_$005 ),
    .set_in_$006    ( areg_file$set_in_$006 ),
    .set_in_$007    ( areg_file$set_in_$007 ),
    .set_in_$008    ( areg_file$set_in_$008 ),
    .set_in_$009    ( areg_file$set_in_$009 ),
    .set_in_$010    ( areg_file$set_in_$010 ),
    .set_in_$011    ( areg_file$set_in_$011 ),
    .set_in_$012    ( areg_file$set_in_$012 ),
    .set_in_$013    ( areg_file$set_in_$013 ),
    .set_in_$014    ( areg_file$set_in_$014 ),
    .set_in_$015    ( areg_file$set_in_$015 ),
    .set_in_$016    ( areg_file$set_in_$016 ),
    .set_in_$017    ( areg_file$set_in_$017 ),
    .set_in_$018    ( areg_file$set_in_$018 ),
    .set_in_$019    ( areg_file$set_in_$019 ),
    .set_in_$020    ( areg_file$set_in_$020 ),
    .set_in_$021    ( areg_file$set_in_$021 ),
    .set_in_$022    ( areg_file$set_in_$022 ),
    .set_in_$023    ( areg_file$set_in_$023 ),
    .set_in_$024    ( areg_file$set_in_$024 ),
    .set_in_$025    ( areg_file$set_in_$025 ),
    .set_in_$026    ( areg_file$set_in_$026 ),
    .set_in_$027    ( areg_file$set_in_$027 ),
    .set_in_$028    ( areg_file$set_in_$028 ),
    .set_in_$029    ( areg_file$set_in_$029 ),
    .set_in_$030    ( areg_file$set_in_$030 ),
    .set_in_$031    ( areg_file$set_in_$031 ),
    .set_call       ( areg_file$set_call ),
    .clk            ( areg_file$clk ),
    .write_addr$000 ( areg_file$write_addr$000 ),
    .read_addr$000  ( areg_file$read_addr$000 ),
    .write_call$000 ( areg_file$write_call$000 ),
    .write_data$000 ( areg_file$write_data$000 ),
    .reset          ( areg_file$reset ),
    .read_data$000  ( areg_file$read_data$000 ),
    .dump_out$000   ( areg_file$dump_out$000 ),
    .dump_out$001   ( areg_file$dump_out$001 ),
    .dump_out$002   ( areg_file$dump_out$002 ),
    .dump_out$003   ( areg_file$dump_out$003 ),
    .dump_out$004   ( areg_file$dump_out$004 ),
    .dump_out$005   ( areg_file$dump_out$005 ),
    .dump_out$006   ( areg_file$dump_out$006 ),
    .dump_out$007   ( areg_file$dump_out$007 ),
    .dump_out$008   ( areg_file$dump_out$008 ),
    .dump_out$009   ( areg_file$dump_out$009 ),
    .dump_out$010   ( areg_file$dump_out$010 ),
    .dump_out$011   ( areg_file$dump_out$011 ),
    .dump_out$012   ( areg_file$dump_out$012 ),
    .dump_out$013   ( areg_file$dump_out$013 ),
    .dump_out$014   ( areg_file$dump_out$014 ),
    .dump_out$015   ( areg_file$dump_out$015 ),
    .dump_out$016   ( areg_file$dump_out$016 ),
    .dump_out$017   ( areg_file$dump_out$017 ),
    .dump_out$018   ( areg_file$dump_out$018 ),
    .dump_out$019   ( areg_file$dump_out$019 ),
    .dump_out$020   ( areg_file$dump_out$020 ),
    .dump_out$021   ( areg_file$dump_out$021 ),
    .dump_out$022   ( areg_file$dump_out$022 ),
    .dump_out$023   ( areg_file$dump_out$023 ),
    .dump_out$024   ( areg_file$dump_out$024 ),
    .dump_out$025   ( areg_file$dump_out$025 ),
    .dump_out$026   ( areg_file$dump_out$026 ),
    .dump_out$027   ( areg_file$dump_out$027 ),
    .dump_out$028   ( areg_file$dump_out$028 ),
    .dump_out$029   ( areg_file$dump_out$029 ),
    .dump_out$030   ( areg_file$dump_out$030 ),
    .dump_out$031   ( areg_file$dump_out$031 )
  );

  // arch_used_pregs temporaries
  logic   [   0:0] arch_used_pregs$set_in_$000;
  logic   [   0:0] arch_used_pregs$set_in_$001;
  logic   [   0:0] arch_used_pregs$set_in_$002;
  logic   [   0:0] arch_used_pregs$set_in_$003;
  logic   [   0:0] arch_used_pregs$set_in_$004;
  logic   [   0:0] arch_used_pregs$set_in_$005;
  logic   [   0:0] arch_used_pregs$set_in_$006;
  logic   [   0:0] arch_used_pregs$set_in_$007;
  logic   [   0:0] arch_used_pregs$set_in_$008;
  logic   [   0:0] arch_used_pregs$set_in_$009;
  logic   [   0:0] arch_used_pregs$set_in_$010;
  logic   [   0:0] arch_used_pregs$set_in_$011;
  logic   [   0:0] arch_used_pregs$set_in_$012;
  logic   [   0:0] arch_used_pregs$set_in_$013;
  logic   [   0:0] arch_used_pregs$set_in_$014;
  logic   [   0:0] arch_used_pregs$set_in_$015;
  logic   [   0:0] arch_used_pregs$set_in_$016;
  logic   [   0:0] arch_used_pregs$set_in_$017;
  logic   [   0:0] arch_used_pregs$set_in_$018;
  logic   [   0:0] arch_used_pregs$set_in_$019;
  logic   [   0:0] arch_used_pregs$set_in_$020;
  logic   [   0:0] arch_used_pregs$set_in_$021;
  logic   [   0:0] arch_used_pregs$set_in_$022;
  logic   [   0:0] arch_used_pregs$set_in_$023;
  logic   [   0:0] arch_used_pregs$set_in_$024;
  logic   [   0:0] arch_used_pregs$set_in_$025;
  logic   [   0:0] arch_used_pregs$set_in_$026;
  logic   [   0:0] arch_used_pregs$set_in_$027;
  logic   [   0:0] arch_used_pregs$set_in_$028;
  logic   [   0:0] arch_used_pregs$set_in_$029;
  logic   [   0:0] arch_used_pregs$set_in_$030;
  logic   [   0:0] arch_used_pregs$set_in_$031;
  logic   [   0:0] arch_used_pregs$set_in_$032;
  logic   [   0:0] arch_used_pregs$set_in_$033;
  logic   [   0:0] arch_used_pregs$set_in_$034;
  logic   [   0:0] arch_used_pregs$set_in_$035;
  logic   [   0:0] arch_used_pregs$set_in_$036;
  logic   [   0:0] arch_used_pregs$set_in_$037;
  logic   [   0:0] arch_used_pregs$set_in_$038;
  logic   [   0:0] arch_used_pregs$set_in_$039;
  logic   [   0:0] arch_used_pregs$set_in_$040;
  logic   [   0:0] arch_used_pregs$set_in_$041;
  logic   [   0:0] arch_used_pregs$set_in_$042;
  logic   [   0:0] arch_used_pregs$set_in_$043;
  logic   [   0:0] arch_used_pregs$set_in_$044;
  logic   [   0:0] arch_used_pregs$set_in_$045;
  logic   [   0:0] arch_used_pregs$set_in_$046;
  logic   [   0:0] arch_used_pregs$set_in_$047;
  logic   [   0:0] arch_used_pregs$set_in_$048;
  logic   [   0:0] arch_used_pregs$set_in_$049;
  logic   [   0:0] arch_used_pregs$set_in_$050;
  logic   [   0:0] arch_used_pregs$set_in_$051;
  logic   [   0:0] arch_used_pregs$set_in_$052;
  logic   [   0:0] arch_used_pregs$set_in_$053;
  logic   [   0:0] arch_used_pregs$set_in_$054;
  logic   [   0:0] arch_used_pregs$set_in_$055;
  logic   [   0:0] arch_used_pregs$set_in_$056;
  logic   [   0:0] arch_used_pregs$set_in_$057;
  logic   [   0:0] arch_used_pregs$set_in_$058;
  logic   [   0:0] arch_used_pregs$set_in_$059;
  logic   [   0:0] arch_used_pregs$set_in_$060;
  logic   [   0:0] arch_used_pregs$set_in_$061;
  logic   [   0:0] arch_used_pregs$set_in_$062;
  logic   [   0:0] arch_used_pregs$set_call;
  logic   [   0:0] arch_used_pregs$clk;
  logic   [   5:0] arch_used_pregs$write_addr$000;
  logic   [   5:0] arch_used_pregs$write_addr$001;
  logic   [   0:0] arch_used_pregs$write_call$000;
  logic   [   0:0] arch_used_pregs$write_call$001;
  logic   [   0:0] arch_used_pregs$write_data$000;
  logic   [   0:0] arch_used_pregs$write_data$001;
  logic   [   0:0] arch_used_pregs$reset;
  logic   [   0:0] arch_used_pregs$dump_out$000;
  logic   [   0:0] arch_used_pregs$dump_out$001;
  logic   [   0:0] arch_used_pregs$dump_out$002;
  logic   [   0:0] arch_used_pregs$dump_out$003;
  logic   [   0:0] arch_used_pregs$dump_out$004;
  logic   [   0:0] arch_used_pregs$dump_out$005;
  logic   [   0:0] arch_used_pregs$dump_out$006;
  logic   [   0:0] arch_used_pregs$dump_out$007;
  logic   [   0:0] arch_used_pregs$dump_out$008;
  logic   [   0:0] arch_used_pregs$dump_out$009;
  logic   [   0:0] arch_used_pregs$dump_out$010;
  logic   [   0:0] arch_used_pregs$dump_out$011;
  logic   [   0:0] arch_used_pregs$dump_out$012;
  logic   [   0:0] arch_used_pregs$dump_out$013;
  logic   [   0:0] arch_used_pregs$dump_out$014;
  logic   [   0:0] arch_used_pregs$dump_out$015;
  logic   [   0:0] arch_used_pregs$dump_out$016;
  logic   [   0:0] arch_used_pregs$dump_out$017;
  logic   [   0:0] arch_used_pregs$dump_out$018;
  logic   [   0:0] arch_used_pregs$dump_out$019;
  logic   [   0:0] arch_used_pregs$dump_out$020;
  logic   [   0:0] arch_used_pregs$dump_out$021;
  logic   [   0:0] arch_used_pregs$dump_out$022;
  logic   [   0:0] arch_used_pregs$dump_out$023;
  logic   [   0:0] arch_used_pregs$dump_out$024;
  logic   [   0:0] arch_used_pregs$dump_out$025;
  logic   [   0:0] arch_used_pregs$dump_out$026;
  logic   [   0:0] arch_used_pregs$dump_out$027;
  logic   [   0:0] arch_used_pregs$dump_out$028;
  logic   [   0:0] arch_used_pregs$dump_out$029;
  logic   [   0:0] arch_used_pregs$dump_out$030;
  logic   [   0:0] arch_used_pregs$dump_out$031;
  logic   [   0:0] arch_used_pregs$dump_out$032;
  logic   [   0:0] arch_used_pregs$dump_out$033;
  logic   [   0:0] arch_used_pregs$dump_out$034;
  logic   [   0:0] arch_used_pregs$dump_out$035;
  logic   [   0:0] arch_used_pregs$dump_out$036;
  logic   [   0:0] arch_used_pregs$dump_out$037;
  logic   [   0:0] arch_used_pregs$dump_out$038;
  logic   [   0:0] arch_used_pregs$dump_out$039;
  logic   [   0:0] arch_used_pregs$dump_out$040;
  logic   [   0:0] arch_used_pregs$dump_out$041;
  logic   [   0:0] arch_used_pregs$dump_out$042;
  logic   [   0:0] arch_used_pregs$dump_out$043;
  logic   [   0:0] arch_used_pregs$dump_out$044;
  logic   [   0:0] arch_used_pregs$dump_out$045;
  logic   [   0:0] arch_used_pregs$dump_out$046;
  logic   [   0:0] arch_used_pregs$dump_out$047;
  logic   [   0:0] arch_used_pregs$dump_out$048;
  logic   [   0:0] arch_used_pregs$dump_out$049;
  logic   [   0:0] arch_used_pregs$dump_out$050;
  logic   [   0:0] arch_used_pregs$dump_out$051;
  logic   [   0:0] arch_used_pregs$dump_out$052;
  logic   [   0:0] arch_used_pregs$dump_out$053;
  logic   [   0:0] arch_used_pregs$dump_out$054;
  logic   [   0:0] arch_used_pregs$dump_out$055;
  logic   [   0:0] arch_used_pregs$dump_out$056;
  logic   [   0:0] arch_used_pregs$dump_out$057;
  logic   [   0:0] arch_used_pregs$dump_out$058;
  logic   [   0:0] arch_used_pregs$dump_out$059;
  logic   [   0:0] arch_used_pregs$dump_out$060;
  logic   [   0:0] arch_used_pregs$dump_out$061;
  logic   [   0:0] arch_used_pregs$dump_out$062;

  RegisterFile_0x39d647b3aea936a6 arch_used_pregs
  (
    .set_in_$000    ( arch_used_pregs$set_in_$000 ),
    .set_in_$001    ( arch_used_pregs$set_in_$001 ),
    .set_in_$002    ( arch_used_pregs$set_in_$002 ),
    .set_in_$003    ( arch_used_pregs$set_in_$003 ),
    .set_in_$004    ( arch_used_pregs$set_in_$004 ),
    .set_in_$005    ( arch_used_pregs$set_in_$005 ),
    .set_in_$006    ( arch_used_pregs$set_in_$006 ),
    .set_in_$007    ( arch_used_pregs$set_in_$007 ),
    .set_in_$008    ( arch_used_pregs$set_in_$008 ),
    .set_in_$009    ( arch_used_pregs$set_in_$009 ),
    .set_in_$010    ( arch_used_pregs$set_in_$010 ),
    .set_in_$011    ( arch_used_pregs$set_in_$011 ),
    .set_in_$012    ( arch_used_pregs$set_in_$012 ),
    .set_in_$013    ( arch_used_pregs$set_in_$013 ),
    .set_in_$014    ( arch_used_pregs$set_in_$014 ),
    .set_in_$015    ( arch_used_pregs$set_in_$015 ),
    .set_in_$016    ( arch_used_pregs$set_in_$016 ),
    .set_in_$017    ( arch_used_pregs$set_in_$017 ),
    .set_in_$018    ( arch_used_pregs$set_in_$018 ),
    .set_in_$019    ( arch_used_pregs$set_in_$019 ),
    .set_in_$020    ( arch_used_pregs$set_in_$020 ),
    .set_in_$021    ( arch_used_pregs$set_in_$021 ),
    .set_in_$022    ( arch_used_pregs$set_in_$022 ),
    .set_in_$023    ( arch_used_pregs$set_in_$023 ),
    .set_in_$024    ( arch_used_pregs$set_in_$024 ),
    .set_in_$025    ( arch_used_pregs$set_in_$025 ),
    .set_in_$026    ( arch_used_pregs$set_in_$026 ),
    .set_in_$027    ( arch_used_pregs$set_in_$027 ),
    .set_in_$028    ( arch_used_pregs$set_in_$028 ),
    .set_in_$029    ( arch_used_pregs$set_in_$029 ),
    .set_in_$030    ( arch_used_pregs$set_in_$030 ),
    .set_in_$031    ( arch_used_pregs$set_in_$031 ),
    .set_in_$032    ( arch_used_pregs$set_in_$032 ),
    .set_in_$033    ( arch_used_pregs$set_in_$033 ),
    .set_in_$034    ( arch_used_pregs$set_in_$034 ),
    .set_in_$035    ( arch_used_pregs$set_in_$035 ),
    .set_in_$036    ( arch_used_pregs$set_in_$036 ),
    .set_in_$037    ( arch_used_pregs$set_in_$037 ),
    .set_in_$038    ( arch_used_pregs$set_in_$038 ),
    .set_in_$039    ( arch_used_pregs$set_in_$039 ),
    .set_in_$040    ( arch_used_pregs$set_in_$040 ),
    .set_in_$041    ( arch_used_pregs$set_in_$041 ),
    .set_in_$042    ( arch_used_pregs$set_in_$042 ),
    .set_in_$043    ( arch_used_pregs$set_in_$043 ),
    .set_in_$044    ( arch_used_pregs$set_in_$044 ),
    .set_in_$045    ( arch_used_pregs$set_in_$045 ),
    .set_in_$046    ( arch_used_pregs$set_in_$046 ),
    .set_in_$047    ( arch_used_pregs$set_in_$047 ),
    .set_in_$048    ( arch_used_pregs$set_in_$048 ),
    .set_in_$049    ( arch_used_pregs$set_in_$049 ),
    .set_in_$050    ( arch_used_pregs$set_in_$050 ),
    .set_in_$051    ( arch_used_pregs$set_in_$051 ),
    .set_in_$052    ( arch_used_pregs$set_in_$052 ),
    .set_in_$053    ( arch_used_pregs$set_in_$053 ),
    .set_in_$054    ( arch_used_pregs$set_in_$054 ),
    .set_in_$055    ( arch_used_pregs$set_in_$055 ),
    .set_in_$056    ( arch_used_pregs$set_in_$056 ),
    .set_in_$057    ( arch_used_pregs$set_in_$057 ),
    .set_in_$058    ( arch_used_pregs$set_in_$058 ),
    .set_in_$059    ( arch_used_pregs$set_in_$059 ),
    .set_in_$060    ( arch_used_pregs$set_in_$060 ),
    .set_in_$061    ( arch_used_pregs$set_in_$061 ),
    .set_in_$062    ( arch_used_pregs$set_in_$062 ),
    .set_call       ( arch_used_pregs$set_call ),
    .clk            ( arch_used_pregs$clk ),
    .write_addr$000 ( arch_used_pregs$write_addr$000 ),
    .write_addr$001 ( arch_used_pregs$write_addr$001 ),
    .write_call$000 ( arch_used_pregs$write_call$000 ),
    .write_call$001 ( arch_used_pregs$write_call$001 ),
    .write_data$000 ( arch_used_pregs$write_data$000 ),
    .write_data$001 ( arch_used_pregs$write_data$001 ),
    .reset          ( arch_used_pregs$reset ),
    .dump_out$000   ( arch_used_pregs$dump_out$000 ),
    .dump_out$001   ( arch_used_pregs$dump_out$001 ),
    .dump_out$002   ( arch_used_pregs$dump_out$002 ),
    .dump_out$003   ( arch_used_pregs$dump_out$003 ),
    .dump_out$004   ( arch_used_pregs$dump_out$004 ),
    .dump_out$005   ( arch_used_pregs$dump_out$005 ),
    .dump_out$006   ( arch_used_pregs$dump_out$006 ),
    .dump_out$007   ( arch_used_pregs$dump_out$007 ),
    .dump_out$008   ( arch_used_pregs$dump_out$008 ),
    .dump_out$009   ( arch_used_pregs$dump_out$009 ),
    .dump_out$010   ( arch_used_pregs$dump_out$010 ),
    .dump_out$011   ( arch_used_pregs$dump_out$011 ),
    .dump_out$012   ( arch_used_pregs$dump_out$012 ),
    .dump_out$013   ( arch_used_pregs$dump_out$013 ),
    .dump_out$014   ( arch_used_pregs$dump_out$014 ),
    .dump_out$015   ( arch_used_pregs$dump_out$015 ),
    .dump_out$016   ( arch_used_pregs$dump_out$016 ),
    .dump_out$017   ( arch_used_pregs$dump_out$017 ),
    .dump_out$018   ( arch_used_pregs$dump_out$018 ),
    .dump_out$019   ( arch_used_pregs$dump_out$019 ),
    .dump_out$020   ( arch_used_pregs$dump_out$020 ),
    .dump_out$021   ( arch_used_pregs$dump_out$021 ),
    .dump_out$022   ( arch_used_pregs$dump_out$022 ),
    .dump_out$023   ( arch_used_pregs$dump_out$023 ),
    .dump_out$024   ( arch_used_pregs$dump_out$024 ),
    .dump_out$025   ( arch_used_pregs$dump_out$025 ),
    .dump_out$026   ( arch_used_pregs$dump_out$026 ),
    .dump_out$027   ( arch_used_pregs$dump_out$027 ),
    .dump_out$028   ( arch_used_pregs$dump_out$028 ),
    .dump_out$029   ( arch_used_pregs$dump_out$029 ),
    .dump_out$030   ( arch_used_pregs$dump_out$030 ),
    .dump_out$031   ( arch_used_pregs$dump_out$031 ),
    .dump_out$032   ( arch_used_pregs$dump_out$032 ),
    .dump_out$033   ( arch_used_pregs$dump_out$033 ),
    .dump_out$034   ( arch_used_pregs$dump_out$034 ),
    .dump_out$035   ( arch_used_pregs$dump_out$035 ),
    .dump_out$036   ( arch_used_pregs$dump_out$036 ),
    .dump_out$037   ( arch_used_pregs$dump_out$037 ),
    .dump_out$038   ( arch_used_pregs$dump_out$038 ),
    .dump_out$039   ( arch_used_pregs$dump_out$039 ),
    .dump_out$040   ( arch_used_pregs$dump_out$040 ),
    .dump_out$041   ( arch_used_pregs$dump_out$041 ),
    .dump_out$042   ( arch_used_pregs$dump_out$042 ),
    .dump_out$043   ( arch_used_pregs$dump_out$043 ),
    .dump_out$044   ( arch_used_pregs$dump_out$044 ),
    .dump_out$045   ( arch_used_pregs$dump_out$045 ),
    .dump_out$046   ( arch_used_pregs$dump_out$046 ),
    .dump_out$047   ( arch_used_pregs$dump_out$047 ),
    .dump_out$048   ( arch_used_pregs$dump_out$048 ),
    .dump_out$049   ( arch_used_pregs$dump_out$049 ),
    .dump_out$050   ( arch_used_pregs$dump_out$050 ),
    .dump_out$051   ( arch_used_pregs$dump_out$051 ),
    .dump_out$052   ( arch_used_pregs$dump_out$052 ),
    .dump_out$053   ( arch_used_pregs$dump_out$053 ),
    .dump_out$054   ( arch_used_pregs$dump_out$054 ),
    .dump_out$055   ( arch_used_pregs$dump_out$055 ),
    .dump_out$056   ( arch_used_pregs$dump_out$056 ),
    .dump_out$057   ( arch_used_pregs$dump_out$057 ),
    .dump_out$058   ( arch_used_pregs$dump_out$058 ),
    .dump_out$059   ( arch_used_pregs$dump_out$059 ),
    .dump_out$060   ( arch_used_pregs$dump_out$060 ),
    .dump_out$061   ( arch_used_pregs$dump_out$061 ),
    .dump_out$062   ( arch_used_pregs$dump_out$062 )
  );

  // read_muxes_value$000 temporaries
  logic   [  63:0] read_muxes_value$000$mux_in_$000;
  logic   [  63:0] read_muxes_value$000$mux_in_$001;
  logic   [   0:0] read_muxes_value$000$clk;
  logic   [   0:0] read_muxes_value$000$reset;
  logic   [   0:0] read_muxes_value$000$mux_select;
  logic   [  63:0] read_muxes_value$000$mux_out;

  Mux_0x1d47079284a028c3 read_muxes_value$000
  (
    .mux_in_$000 ( read_muxes_value$000$mux_in_$000 ),
    .mux_in_$001 ( read_muxes_value$000$mux_in_$001 ),
    .clk         ( read_muxes_value$000$clk ),
    .reset       ( read_muxes_value$000$reset ),
    .mux_select  ( read_muxes_value$000$mux_select ),
    .mux_out     ( read_muxes_value$000$mux_out )
  );

  // read_muxes_value$001 temporaries
  logic   [  63:0] read_muxes_value$001$mux_in_$000;
  logic   [  63:0] read_muxes_value$001$mux_in_$001;
  logic   [   0:0] read_muxes_value$001$clk;
  logic   [   0:0] read_muxes_value$001$reset;
  logic   [   0:0] read_muxes_value$001$mux_select;
  logic   [  63:0] read_muxes_value$001$mux_out;

  Mux_0x1d47079284a028c3 read_muxes_value$001
  (
    .mux_in_$000 ( read_muxes_value$001$mux_in_$000 ),
    .mux_in_$001 ( read_muxes_value$001$mux_in_$001 ),
    .clk         ( read_muxes_value$001$clk ),
    .reset       ( read_muxes_value$001$reset ),
    .mux_select  ( read_muxes_value$001$mux_select ),
    .mux_out     ( read_muxes_value$001$mux_out )
  );

  // preg_file temporaries
  logic   [   0:0] preg_file$clk;
  logic   [   5:0] preg_file$write_addr$000;
  logic   [   5:0] preg_file$write_addr$001;
  logic   [   5:0] preg_file$read_addr$000;
  logic   [   5:0] preg_file$read_addr$001;
  logic   [   0:0] preg_file$write_call$000;
  logic   [   0:0] preg_file$write_call$001;
  logic   [  63:0] preg_file$write_data$000;
  logic   [  63:0] preg_file$write_data$001;
  logic   [   0:0] preg_file$reset;
  logic   [  63:0] preg_file$read_data$000;
  logic   [  63:0] preg_file$read_data$001;

  AsynchronousRAM_0xb915281a52f5e7 preg_file
  (
    .clk            ( preg_file$clk ),
    .write_addr$000 ( preg_file$write_addr$000 ),
    .write_addr$001 ( preg_file$write_addr$001 ),
    .read_addr$000  ( preg_file$read_addr$000 ),
    .read_addr$001  ( preg_file$read_addr$001 ),
    .write_call$000 ( preg_file$write_call$000 ),
    .write_call$001 ( preg_file$write_call$001 ),
    .write_data$000 ( preg_file$write_data$000 ),
    .write_data$001 ( preg_file$write_data$001 ),
    .reset          ( preg_file$reset ),
    .read_data$000  ( preg_file$read_data$000 ),
    .read_data$001  ( preg_file$read_data$001 )
  );

  // free_regs temporaries
  logic   [   0:0] free_regs$revert_allocs_call;
  logic   [   0:0] free_regs$set_call;
  logic   [   0:0] free_regs$revert_allocs_source_id;
  logic   [   0:0] free_regs$clk;
  logic   [   0:0] free_regs$free_call$000;
  logic   [   0:0] free_regs$free_call$001;
  logic   [   0:0] free_regs$reset_alloc_tracking_call;
  logic   [   0:0] free_regs$reset_alloc_tracking_target_id;
  logic   [   0:0] free_regs$alloc_call$000;
  logic   [   0:0] free_regs$reset;
  logic   [   5:0] free_regs$free_index$000;
  logic   [   5:0] free_regs$free_index$001;
  logic   [  62:0] free_regs$alloc_mask$000;
  logic   [   0:0] free_regs$alloc_rdy$000;
  logic   [   5:0] free_regs$alloc_index$000;

  SnapshottingFreeList_0x68f914e32e2c4f6d free_regs
  (
    .set_state                      ( free_regs$set_state ),
    .revert_allocs_call             ( free_regs$revert_allocs_call ),
    .set_call                       ( free_regs$set_call ),
    .revert_allocs_source_id        ( free_regs$revert_allocs_source_id ),
    .clk                            ( free_regs$clk ),
    .free_call$000                  ( free_regs$free_call$000 ),
    .free_call$001                  ( free_regs$free_call$001 ),
    .reset_alloc_tracking_call      ( free_regs$reset_alloc_tracking_call ),
    .reset_alloc_tracking_target_id ( free_regs$reset_alloc_tracking_target_id ),
    .alloc_call$000                 ( free_regs$alloc_call$000 ),
    .reset                          ( free_regs$reset ),
    .free_index$000                 ( free_regs$free_index$000 ),
    .free_index$001                 ( free_regs$free_index$001 ),
    .alloc_mask$000                 ( free_regs$alloc_mask$000 ),
    .alloc_rdy$000                  ( free_regs$alloc_rdy$000 ),
    .alloc_index$000                ( free_regs$alloc_index$000 )
  );

  // signal connections
  assign arch_used_pregs$clk                               = clk;
  assign arch_used_pregs$reset                             = reset;
  assign arch_used_pregs$write_addr$000                    = areg_file$read_data$000;
  assign arch_used_pregs$write_addr$001                    = commit_tag$000;
  assign arch_used_pregs$write_call$000                    = is_commit_not_zero_tag$000;
  assign arch_used_pregs$write_call$001                    = is_commit_not_zero_tag$000;
  assign arch_used_pregs$write_data$000                    = 1'd0;
  assign arch_used_pregs$write_data$001                    = 1'd1;
  assign arch_used_pregs_packer$clk                        = clk;
  assign arch_used_pregs_packer$pack_in_$000               = arch_used_pregs$dump_out$000;
  assign arch_used_pregs_packer$pack_in_$001               = arch_used_pregs$dump_out$001;
  assign arch_used_pregs_packer$pack_in_$002               = arch_used_pregs$dump_out$002;
  assign arch_used_pregs_packer$pack_in_$003               = arch_used_pregs$dump_out$003;
  assign arch_used_pregs_packer$pack_in_$004               = arch_used_pregs$dump_out$004;
  assign arch_used_pregs_packer$pack_in_$005               = arch_used_pregs$dump_out$005;
  assign arch_used_pregs_packer$pack_in_$006               = arch_used_pregs$dump_out$006;
  assign arch_used_pregs_packer$pack_in_$007               = arch_used_pregs$dump_out$007;
  assign arch_used_pregs_packer$pack_in_$008               = arch_used_pregs$dump_out$008;
  assign arch_used_pregs_packer$pack_in_$009               = arch_used_pregs$dump_out$009;
  assign arch_used_pregs_packer$pack_in_$010               = arch_used_pregs$dump_out$010;
  assign arch_used_pregs_packer$pack_in_$011               = arch_used_pregs$dump_out$011;
  assign arch_used_pregs_packer$pack_in_$012               = arch_used_pregs$dump_out$012;
  assign arch_used_pregs_packer$pack_in_$013               = arch_used_pregs$dump_out$013;
  assign arch_used_pregs_packer$pack_in_$014               = arch_used_pregs$dump_out$014;
  assign arch_used_pregs_packer$pack_in_$015               = arch_used_pregs$dump_out$015;
  assign arch_used_pregs_packer$pack_in_$016               = arch_used_pregs$dump_out$016;
  assign arch_used_pregs_packer$pack_in_$017               = arch_used_pregs$dump_out$017;
  assign arch_used_pregs_packer$pack_in_$018               = arch_used_pregs$dump_out$018;
  assign arch_used_pregs_packer$pack_in_$019               = arch_used_pregs$dump_out$019;
  assign arch_used_pregs_packer$pack_in_$020               = arch_used_pregs$dump_out$020;
  assign arch_used_pregs_packer$pack_in_$021               = arch_used_pregs$dump_out$021;
  assign arch_used_pregs_packer$pack_in_$022               = arch_used_pregs$dump_out$022;
  assign arch_used_pregs_packer$pack_in_$023               = arch_used_pregs$dump_out$023;
  assign arch_used_pregs_packer$pack_in_$024               = arch_used_pregs$dump_out$024;
  assign arch_used_pregs_packer$pack_in_$025               = arch_used_pregs$dump_out$025;
  assign arch_used_pregs_packer$pack_in_$026               = arch_used_pregs$dump_out$026;
  assign arch_used_pregs_packer$pack_in_$027               = arch_used_pregs$dump_out$027;
  assign arch_used_pregs_packer$pack_in_$028               = arch_used_pregs$dump_out$028;
  assign arch_used_pregs_packer$pack_in_$029               = arch_used_pregs$dump_out$029;
  assign arch_used_pregs_packer$pack_in_$030               = arch_used_pregs$dump_out$030;
  assign arch_used_pregs_packer$pack_in_$031               = arch_used_pregs$dump_out$031;
  assign arch_used_pregs_packer$pack_in_$032               = arch_used_pregs$dump_out$032;
  assign arch_used_pregs_packer$pack_in_$033               = arch_used_pregs$dump_out$033;
  assign arch_used_pregs_packer$pack_in_$034               = arch_used_pregs$dump_out$034;
  assign arch_used_pregs_packer$pack_in_$035               = arch_used_pregs$dump_out$035;
  assign arch_used_pregs_packer$pack_in_$036               = arch_used_pregs$dump_out$036;
  assign arch_used_pregs_packer$pack_in_$037               = arch_used_pregs$dump_out$037;
  assign arch_used_pregs_packer$pack_in_$038               = arch_used_pregs$dump_out$038;
  assign arch_used_pregs_packer$pack_in_$039               = arch_used_pregs$dump_out$039;
  assign arch_used_pregs_packer$pack_in_$040               = arch_used_pregs$dump_out$040;
  assign arch_used_pregs_packer$pack_in_$041               = arch_used_pregs$dump_out$041;
  assign arch_used_pregs_packer$pack_in_$042               = arch_used_pregs$dump_out$042;
  assign arch_used_pregs_packer$pack_in_$043               = arch_used_pregs$dump_out$043;
  assign arch_used_pregs_packer$pack_in_$044               = arch_used_pregs$dump_out$044;
  assign arch_used_pregs_packer$pack_in_$045               = arch_used_pregs$dump_out$045;
  assign arch_used_pregs_packer$pack_in_$046               = arch_used_pregs$dump_out$046;
  assign arch_used_pregs_packer$pack_in_$047               = arch_used_pregs$dump_out$047;
  assign arch_used_pregs_packer$pack_in_$048               = arch_used_pregs$dump_out$048;
  assign arch_used_pregs_packer$pack_in_$049               = arch_used_pregs$dump_out$049;
  assign arch_used_pregs_packer$pack_in_$050               = arch_used_pregs$dump_out$050;
  assign arch_used_pregs_packer$pack_in_$051               = arch_used_pregs$dump_out$051;
  assign arch_used_pregs_packer$pack_in_$052               = arch_used_pregs$dump_out$052;
  assign arch_used_pregs_packer$pack_in_$053               = arch_used_pregs$dump_out$053;
  assign arch_used_pregs_packer$pack_in_$054               = arch_used_pregs$dump_out$054;
  assign arch_used_pregs_packer$pack_in_$055               = arch_used_pregs$dump_out$055;
  assign arch_used_pregs_packer$pack_in_$056               = arch_used_pregs$dump_out$056;
  assign arch_used_pregs_packer$pack_in_$057               = arch_used_pregs$dump_out$057;
  assign arch_used_pregs_packer$pack_in_$058               = arch_used_pregs$dump_out$058;
  assign arch_used_pregs_packer$pack_in_$059               = arch_used_pregs$dump_out$059;
  assign arch_used_pregs_packer$pack_in_$060               = arch_used_pregs$dump_out$060;
  assign arch_used_pregs_packer$pack_in_$061               = arch_used_pregs$dump_out$061;
  assign arch_used_pregs_packer$pack_in_$062               = arch_used_pregs$dump_out$062;
  assign arch_used_pregs_packer$reset                      = reset;
  assign areg_file$clk                                     = clk;
  assign areg_file$read_addr$000                           = inverse$read_data$000;
  assign areg_file$reset                                   = reset;
  assign areg_file$write_addr$000                          = inverse$read_data$000;
  assign areg_file$write_call$000                          = is_commit_not_zero_tag$000;
  assign areg_file$write_data$000                          = commit_tag$000;
  assign free_regs$clk                                     = clk;
  assign free_regs$free_call$000                           = is_commit_not_zero_tag$000;
  assign free_regs$free_index$000                          = areg_file$read_data$000;
  assign free_regs$reset                                   = reset;
  assign free_regs$reset_alloc_tracking_call               = snapshot_call;
  assign free_regs$reset_alloc_tracking_target_id          = snapshot_id_;
  assign free_regs$revert_allocs_call                      = restore_call;
  assign free_regs$revert_allocs_source_id                 = restore_source_id;
  assign free_regs$set_call                                = rollback_call;
  assign get_dst_rdy$000                                   = free_regs$alloc_rdy$000;
  assign get_src_preg$000                                  = rename_table$lookup_preg$000;
  assign get_src_preg$001                                  = rename_table$lookup_preg$001;
  assign get_updated_incremental_masks$000                 = 64'd0;
  assign get_updated_mask                                  = get_updated_incremental_masks$001;
  assign inverse$clk                                       = clk;
  assign inverse$read_addr$000                             = commit_tag$000;
  assign inverse$reset                                     = reset;
  assign inverse$write_addr$000                            = get_dst_preg$000;
  assign inverse$write_call$000                            = get_dst_need_writeback$000;
  assign inverse$write_data$000                            = get_dst_areg$000;
  assign is_ready_ready$000                                = read_muxes_ready$000$mux_out;
  assign is_ready_ready$001                                = read_muxes_ready$001$mux_out;
  assign preg_file$clk                                     = clk;
  assign preg_file$read_addr$000                           = read_tag$000;
  assign preg_file$read_addr$001                           = read_tag$001;
  assign preg_file$reset                                   = reset;
  assign preg_file$write_addr$000                          = write_tag$000;
  assign preg_file$write_addr$001                          = get_dst_preg$000;
  assign preg_file$write_call$000                          = is_write_not_zero_tag$000;
  assign preg_file$write_call$001                          = get_dst_need_writeback$000;
  assign preg_file$write_data$000                          = write_value$000;
  assign preg_file$write_data$001                          = 64'd0;
  assign read_muxes_ready$000$clk                          = clk;
  assign read_muxes_ready$000$mux_in_$000                  = ready_table$read_data$000;
  assign read_muxes_ready$000$mux_in_$001                  = 1'd1;
  assign read_muxes_ready$000$mux_select                   = is_ready_is_zero_tag$000;
  assign read_muxes_ready$000$reset                        = reset;
  assign read_muxes_ready$001$clk                          = clk;
  assign read_muxes_ready$001$mux_in_$000                  = ready_table$read_data$001;
  assign read_muxes_ready$001$mux_in_$001                  = 1'd1;
  assign read_muxes_ready$001$mux_select                   = is_ready_is_zero_tag$001;
  assign read_muxes_ready$001$reset                        = reset;
  assign read_muxes_value$000$clk                          = clk;
  assign read_muxes_value$000$mux_in_$000                  = preg_file$read_data$000;
  assign read_muxes_value$000$mux_in_$001                  = 64'd0;
  assign read_muxes_value$000$mux_select                   = read_is_zero_tag$000;
  assign read_muxes_value$000$reset                        = reset;
  assign read_muxes_value$001$clk                          = clk;
  assign read_muxes_value$001$mux_in_$000                  = preg_file$read_data$001;
  assign read_muxes_value$001$mux_in_$001                  = 64'd0;
  assign read_muxes_value$001$mux_select                   = read_is_zero_tag$001;
  assign read_muxes_value$001$reset                        = reset;
  assign read_value$000                                    = read_muxes_value$000$mux_out;
  assign read_value$001                                    = read_muxes_value$001$mux_out;
  assign ready_table$clk                                   = clk;
  assign ready_table$read_addr$000                         = is_ready_tag$000;
  assign ready_table$read_addr$001                         = is_ready_tag$001;
  assign ready_table$reset                                 = reset;
  assign ready_table$write_addr$000                        = write_tag$000;
  assign ready_table$write_addr$001                        = get_dst_preg$000;
  assign ready_table$write_call$000                        = is_write_not_zero_tag$000;
  assign ready_table$write_call$001                        = get_dst_need_writeback$000;
  assign ready_table$write_data$000                        = 1'd1;
  assign ready_table$write_data$001                        = 1'd0;
  assign rename_table$clk                                  = clk;
  assign rename_table$lookup_areg$000                      = get_src_areg$000;
  assign rename_table$lookup_areg$001                      = get_src_areg$001;
  assign rename_table$reset                                = reset;
  assign rename_table$restore_call                         = restore_call;
  assign rename_table$restore_source_id                    = restore_source_id;
  assign rename_table$set_call                             = rollback_call;
  assign rename_table$set_in_$000                          = areg_file$dump_out$000;
  assign rename_table$set_in_$001                          = areg_file$dump_out$001;
  assign rename_table$set_in_$002                          = areg_file$dump_out$002;
  assign rename_table$set_in_$003                          = areg_file$dump_out$003;
  assign rename_table$set_in_$004                          = areg_file$dump_out$004;
  assign rename_table$set_in_$005                          = areg_file$dump_out$005;
  assign rename_table$set_in_$006                          = areg_file$dump_out$006;
  assign rename_table$set_in_$007                          = areg_file$dump_out$007;
  assign rename_table$set_in_$008                          = areg_file$dump_out$008;
  assign rename_table$set_in_$009                          = areg_file$dump_out$009;
  assign rename_table$set_in_$010                          = areg_file$dump_out$010;
  assign rename_table$set_in_$011                          = areg_file$dump_out$011;
  assign rename_table$set_in_$012                          = areg_file$dump_out$012;
  assign rename_table$set_in_$013                          = areg_file$dump_out$013;
  assign rename_table$set_in_$014                          = areg_file$dump_out$014;
  assign rename_table$set_in_$015                          = areg_file$dump_out$015;
  assign rename_table$set_in_$016                          = areg_file$dump_out$016;
  assign rename_table$set_in_$017                          = areg_file$dump_out$017;
  assign rename_table$set_in_$018                          = areg_file$dump_out$018;
  assign rename_table$set_in_$019                          = areg_file$dump_out$019;
  assign rename_table$set_in_$020                          = areg_file$dump_out$020;
  assign rename_table$set_in_$021                          = areg_file$dump_out$021;
  assign rename_table$set_in_$022                          = areg_file$dump_out$022;
  assign rename_table$set_in_$023                          = areg_file$dump_out$023;
  assign rename_table$set_in_$024                          = areg_file$dump_out$024;
  assign rename_table$set_in_$025                          = areg_file$dump_out$025;
  assign rename_table$set_in_$026                          = areg_file$dump_out$026;
  assign rename_table$set_in_$027                          = areg_file$dump_out$027;
  assign rename_table$set_in_$028                          = areg_file$dump_out$028;
  assign rename_table$set_in_$029                          = areg_file$dump_out$029;
  assign rename_table$set_in_$030                          = areg_file$dump_out$030;
  assign rename_table$set_in_$031                          = areg_file$dump_out$031;
  assign rename_table$snapshot_call                        = snapshot_call;
  assign rename_table$snapshot_target_id                   = snapshot_id_;
  assign rename_table$update_areg$000                      = get_dst_areg$000;
  assign rename_table$update_call$000                      = get_dst_need_writeback$000;
  assign rename_table$update_preg$000                      = get_dst_preg$000;
  assign snapshot_allocator$alloc_call$000                 = snapshot_call;
  assign snapshot_allocator$clk                            = clk;
  assign snapshot_allocator$free_call$000                  = free_snapshot_call;
  assign snapshot_allocator$free_index$000                 = free_snapshot_id_;
  assign snapshot_allocator$reset                          = reset;
  assign snapshot_allocator$reset_alloc_tracking_call      = snapshot_call;
  assign snapshot_allocator$reset_alloc_tracking_target_id = snapshot_id_;
  assign snapshot_allocator$revert_allocs_call             = restore_call;
  assign snapshot_allocator$revert_allocs_source_id        = restore_source_id;
  assign snapshot_allocator$set_call                       = rollback_call;
  assign snapshot_allocator$set_state                      = 2'd3;
  assign snapshot_id_                                      = snapshot_allocator$alloc_index$000;
  assign snapshot_rdy                                      = snapshot_allocator$alloc_rdy$000;

  // array declarations
  logic   [   0:0] commit_call[0:0];
  assign commit_call[  0] = commit_call$000;
  logic   [   5:0] commit_tag[0:0];
  assign commit_tag[  0] = commit_tag$000;
  logic    [   0:0] free_regs$alloc_call[0:0];
  assign free_regs$alloc_call$000 = free_regs$alloc_call[  0];
  logic   [   5:0] free_regs$alloc_index[0:0];
  assign free_regs$alloc_index[  0] = free_regs$alloc_index$000;
  logic   [   0:0] free_regs$alloc_rdy[0:0];
  assign free_regs$alloc_rdy[  0] = free_regs$alloc_rdy$000;
  logic   [   4:0] get_dst_areg[0:0];
  assign get_dst_areg[  0] = get_dst_areg$000;
  logic   [   0:0] get_dst_call[0:0];
  assign get_dst_call[  0] = get_dst_call$000;
  logic    [   0:0] get_dst_need_writeback[0:0];
  assign get_dst_need_writeback$000 = get_dst_need_writeback[  0];
  logic    [   5:0] get_dst_preg[0:0];
  assign get_dst_preg$000 = get_dst_preg[  0];
  logic    [  63:0] get_updated_incremental_masks[0:1];
  assign get_updated_incremental_masks$000 = get_updated_incremental_masks[  0];
  assign get_updated_incremental_masks$001 = get_updated_incremental_masks[  1];
  logic    [   0:0] is_commit_not_zero_tag[0:0];
  assign is_commit_not_zero_tag$000 = is_commit_not_zero_tag[  0];
  logic    [   0:0] is_ready_is_zero_tag[0:1];
  assign is_ready_is_zero_tag$000 = is_ready_is_zero_tag[  0];
  assign is_ready_is_zero_tag$001 = is_ready_is_zero_tag[  1];
  logic   [   5:0] is_ready_tag[0:1];
  assign is_ready_tag[  0] = is_ready_tag$000;
  assign is_ready_tag[  1] = is_ready_tag$001;
  logic    [   0:0] is_write_not_zero_tag[0:0];
  assign is_write_not_zero_tag$000 = is_write_not_zero_tag[  0];
  logic    [   0:0] read_is_zero_tag[0:1];
  assign read_is_zero_tag$000 = read_is_zero_tag[  0];
  assign read_is_zero_tag$001 = read_is_zero_tag[  1];
  logic   [   5:0] read_tag[0:1];
  assign read_tag[  0] = read_tag$000;
  assign read_tag[  1] = read_tag$001;
  logic   [   0:0] write_call[0:0];
  assign write_call[  0] = write_call$000;
  logic   [   5:0] write_tag[0:0];
  assign write_tag[  0] = write_tag$000;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def check_commit(i=i):
  //         s.is_commit_not_zero_tag[i].v = (s.commit_tag[i] !=
  //                                          s.ZERO_TAG) and s.commit_call[i]

  // logic for check_commit()
  always @ (*) begin
    is_commit_not_zero_tag[0] = ((commit_tag[0] != ZERO_TAG)&&commit_call[0]);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def check_write(i=i):
  //         s.is_write_not_zero_tag[i].v = (s.write_tag[i] !=
  //                                         s.ZERO_TAG) and s.write_call[i]

  // logic for check_write()
  always @ (*) begin
    is_write_not_zero_tag[0] = ((write_tag[0] != ZERO_TAG)&&write_call[0]);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def get_updated_mask(curr=i + 1, last=i):
  //         s.get_updated_incremental_masks[
  //             curr].v = s.get_updated_incremental_masks[last]
  //         if s.is_write_not_zero_tag[last]:
  //           s.get_updated_incremental_masks[curr][s.write_tag[last]].v = 1

  // logic for get_updated_mask()
  always @ (*) begin
    get_updated_incremental_masks[1] = get_updated_incremental_masks[0];
    if (is_write_not_zero_tag[0]) begin
      get_updated_incremental_masks[1][write_tag[0]] = 1;
    end
    else begin
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_get_dst_allocate(i=i):
  //         if s.get_dst_areg[i] == 0:
  //           # zero register
  //           s.free_regs.alloc_call[i].v = 0
  //           s.get_dst_preg[i].v = s.ZERO_TAG
  //           s.get_dst_need_writeback[i].v = 0
  //         elif s.free_regs.alloc_rdy[i]:
  //           # allocate a register from the freelist
  //           s.free_regs.alloc_call[i].v = s.get_dst_call[i]
  //           s.get_dst_preg[i].v = s.free_regs.alloc_index[i]
  //           s.get_dst_need_writeback[i].v = s.get_dst_call[i]
  //         else:
  //           # free list is full
  //           s.free_regs.alloc_call[i].v = 0
  //           s.get_dst_preg[i].v = s.ZERO_TAG
  //           s.get_dst_need_writeback[i].v = 0

  // logic for handle_get_dst_allocate()
  always @ (*) begin
    if ((get_dst_areg[0] == 0)) begin
      free_regs$alloc_call[0] = 0;
      get_dst_preg[0] = ZERO_TAG;
      get_dst_need_writeback[0] = 0;
    end
    else begin
      if (free_regs$alloc_rdy[0]) begin
        free_regs$alloc_call[0] = get_dst_call[0];
        get_dst_preg[0] = free_regs$alloc_index[0];
        get_dst_need_writeback[0] = get_dst_call[0];
      end
      else begin
        free_regs$alloc_call[0] = 0;
        get_dst_preg[0] = ZERO_TAG;
        get_dst_need_writeback[0] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_read(i=i):
  //         s.is_ready_is_zero_tag[i].v = s.is_ready_tag[i] == s.ZERO_TAG

  // logic for handle_read()
  always @ (*) begin
    is_ready_is_zero_tag[0] = (is_ready_tag[0] == ZERO_TAG);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_read(i=i):
  //         s.is_ready_is_zero_tag[i].v = s.is_ready_tag[i] == s.ZERO_TAG

  // logic for handle_read()
  always @ (*) begin
    is_ready_is_zero_tag[1] = (is_ready_tag[1] == ZERO_TAG);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_read(i=i):
  //         s.read_is_zero_tag[i].v = s.read_tag[i] == s.ZERO_TAG

  // logic for handle_read()
  always @ (*) begin
    read_is_zero_tag[0] = (read_tag[0] == ZERO_TAG);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_read(i=i):
  //         s.read_is_zero_tag[i].v = s.read_tag[i] == s.ZERO_TAG

  // logic for handle_read()
  always @ (*) begin
    read_is_zero_tag[1] = (read_tag[1] == ZERO_TAG);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_rollback_free_regs_set():
  //       s.free_regs.set_state.v = ~s.arch_used_pregs_packer.pack_packed

  // logic for handle_rollback_free_regs_set()
  always @ (*) begin
    free_regs$set_state = ~arch_used_pregs_packer$pack_packed;
  end


endmodule // DataFlowManager_0x54912d9190dab9c9

//-----------------------------------------------------------------------------
// SnapshottingFreeList_0x64ee202bb6767a5b
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.snapshotting_freelist {"freelist_impl": "<class 'util.rtl.freelist.FreeList'>", "nslots": 2, "nsnapshots": 2, "num_alloc_ports": 1, "num_free_ports": 1, "used_slots_initial": 0}
// PyMTL: verilator_xinit = zeros
module SnapshottingFreeList_0x64ee202bb6767a5b
(
  input  logic [   0:0] alloc_call$000,
  output logic [   0:0] alloc_index$000,
  output logic [   1:0] alloc_mask$000,
  output logic [   0:0] alloc_rdy$000,
  input  logic [   0:0] clk,
  input  logic [   0:0] free_call$000,
  input  logic [   0:0] free_index$000,
  input  logic [   0:0] reset,
  input  logic [   0:0] reset_alloc_tracking_call,
  input  logic [   0:0] reset_alloc_tracking_target_id,
  input  logic [   0:0] revert_allocs_call,
  input  logic [   0:0] revert_allocs_source_id,
  input  logic [   0:0] set_call,
  input  logic [   1:0] set_state
);

  // register declarations
  logic    [   0:0] free_list$release_call;

  // snapshots$000 temporaries
  logic   [   0:0] snapshots$000$set_in_$000;
  logic   [   0:0] snapshots$000$set_in_$001;
  logic   [   0:0] snapshots$000$set_call;
  logic   [   0:0] snapshots$000$clk;
  logic   [   0:0] snapshots$000$write_addr$000;
  logic   [   0:0] snapshots$000$write_call$000;
  logic   [   0:0] snapshots$000$write_data$000;
  logic   [   0:0] snapshots$000$reset;
  logic   [   0:0] snapshots$000$dump_out$000;
  logic   [   0:0] snapshots$000$dump_out$001;

  RegisterFile_0x6d9ba9c872129f4f snapshots$000
  (
    .set_in_$000    ( snapshots$000$set_in_$000 ),
    .set_in_$001    ( snapshots$000$set_in_$001 ),
    .set_call       ( snapshots$000$set_call ),
    .clk            ( snapshots$000$clk ),
    .write_addr$000 ( snapshots$000$write_addr$000 ),
    .write_call$000 ( snapshots$000$write_call$000 ),
    .write_data$000 ( snapshots$000$write_data$000 ),
    .reset          ( snapshots$000$reset ),
    .dump_out$000   ( snapshots$000$dump_out$000 ),
    .dump_out$001   ( snapshots$000$dump_out$001 )
  );

  // snapshots$001 temporaries
  logic   [   0:0] snapshots$001$set_in_$000;
  logic   [   0:0] snapshots$001$set_in_$001;
  logic   [   0:0] snapshots$001$set_call;
  logic   [   0:0] snapshots$001$clk;
  logic   [   0:0] snapshots$001$write_addr$000;
  logic   [   0:0] snapshots$001$write_call$000;
  logic   [   0:0] snapshots$001$write_data$000;
  logic   [   0:0] snapshots$001$reset;
  logic   [   0:0] snapshots$001$dump_out$000;
  logic   [   0:0] snapshots$001$dump_out$001;

  RegisterFile_0x6d9ba9c872129f4f snapshots$001
  (
    .set_in_$000    ( snapshots$001$set_in_$000 ),
    .set_in_$001    ( snapshots$001$set_in_$001 ),
    .set_call       ( snapshots$001$set_call ),
    .clk            ( snapshots$001$clk ),
    .write_addr$000 ( snapshots$001$write_addr$000 ),
    .write_call$000 ( snapshots$001$write_call$000 ),
    .write_data$000 ( snapshots$001$write_data$000 ),
    .reset          ( snapshots$001$reset ),
    .dump_out$000   ( snapshots$001$dump_out$000 ),
    .dump_out$001   ( snapshots$001$dump_out$001 )
  );

  // dump_mux temporaries
  logic   [   1:0] dump_mux$mux_in_$000;
  logic   [   1:0] dump_mux$mux_in_$001;
  logic   [   0:0] dump_mux$clk;
  logic   [   0:0] dump_mux$reset;
  logic   [   0:0] dump_mux$mux_select;
  logic   [   1:0] dump_mux$mux_out;

  Mux_0x7cc3cbcc1953dfea dump_mux
  (
    .mux_in_$000 ( dump_mux$mux_in_$000 ),
    .mux_in_$001 ( dump_mux$mux_in_$001 ),
    .clk         ( dump_mux$clk ),
    .reset       ( dump_mux$reset ),
    .mux_select  ( dump_mux$mux_select ),
    .mux_out     ( dump_mux$mux_out )
  );

  // free_list temporaries
  logic   [   1:0] free_list$set_state;
  logic   [   0:0] free_list$clk;
  logic   [   0:0] free_list$free_call$000;
  logic   [   1:0] free_list$release_mask;
  logic   [   0:0] free_list$alloc_call$000;
  logic   [   0:0] free_list$reset;
  logic   [   0:0] free_list$set_call;
  logic   [   0:0] free_list$free_index$000;
  logic   [   1:0] free_list$alloc_mask$000;
  logic   [   0:0] free_list$alloc_rdy$000;
  logic   [   0:0] free_list$alloc_index$000;

  FreeList_0x260f6d53b9562731 free_list
  (
    .set_state       ( free_list$set_state ),
    .release_call    ( free_list$release_call ),
    .clk             ( free_list$clk ),
    .free_call$000   ( free_list$free_call$000 ),
    .release_mask    ( free_list$release_mask ),
    .alloc_call$000  ( free_list$alloc_call$000 ),
    .reset           ( free_list$reset ),
    .set_call        ( free_list$set_call ),
    .free_index$000  ( free_list$free_index$000 ),
    .alloc_mask$000  ( free_list$alloc_mask$000 ),
    .alloc_rdy$000   ( free_list$alloc_rdy$000 ),
    .alloc_index$000 ( free_list$alloc_index$000 )
  );

  // snapshot_packers$000 temporaries
  logic   [   0:0] snapshot_packers$000$clk;
  logic   [   0:0] snapshot_packers$000$pack_in_$000;
  logic   [   0:0] snapshot_packers$000$pack_in_$001;
  logic   [   0:0] snapshot_packers$000$reset;
  logic   [   1:0] snapshot_packers$000$pack_packed;

  Packer_0x67209f7520cf166 snapshot_packers$000
  (
    .clk          ( snapshot_packers$000$clk ),
    .pack_in_$000 ( snapshot_packers$000$pack_in_$000 ),
    .pack_in_$001 ( snapshot_packers$000$pack_in_$001 ),
    .reset        ( snapshot_packers$000$reset ),
    .pack_packed  ( snapshot_packers$000$pack_packed )
  );

  // snapshot_packers$001 temporaries
  logic   [   0:0] snapshot_packers$001$clk;
  logic   [   0:0] snapshot_packers$001$pack_in_$000;
  logic   [   0:0] snapshot_packers$001$pack_in_$001;
  logic   [   0:0] snapshot_packers$001$reset;
  logic   [   1:0] snapshot_packers$001$pack_packed;

  Packer_0x67209f7520cf166 snapshot_packers$001
  (
    .clk          ( snapshot_packers$001$clk ),
    .pack_in_$000 ( snapshot_packers$001$pack_in_$000 ),
    .pack_in_$001 ( snapshot_packers$001$pack_in_$001 ),
    .reset        ( snapshot_packers$001$reset ),
    .pack_packed  ( snapshot_packers$001$pack_packed )
  );

  // clean_mux temporaries
  logic   [   1:0] clean_mux$mux_in_$000;
  logic   [   1:0] clean_mux$mux_in_$001;
  logic   [   0:0] clean_mux$clk;
  logic   [   0:0] clean_mux$reset;
  logic   [   0:0] clean_mux$mux_select;
  logic   [   1:0] clean_mux$mux_out;

  Mux_0x7cc3cbcc1953dfea clean_mux
  (
    .mux_in_$000 ( clean_mux$mux_in_$000 ),
    .mux_in_$001 ( clean_mux$mux_in_$001 ),
    .clk         ( clean_mux$clk ),
    .reset       ( clean_mux$reset ),
    .mux_select  ( clean_mux$mux_select ),
    .mux_out     ( clean_mux$mux_out )
  );

  // signal connections
  assign alloc_index$000                   = free_list$alloc_index$000;
  assign alloc_mask$000                    = free_list$alloc_mask$000;
  assign alloc_rdy$000                     = free_list$alloc_rdy$000;
  assign clean_mux$clk                     = clk;
  assign clean_mux$reset                   = reset;
  assign dump_mux$clk                      = clk;
  assign dump_mux$mux_in_$000              = snapshot_packers$000$pack_packed;
  assign dump_mux$mux_in_$001              = snapshot_packers$001$pack_packed;
  assign dump_mux$mux_select               = revert_allocs_source_id;
  assign dump_mux$reset                    = reset;
  assign free_list$alloc_call$000          = alloc_call$000;
  assign free_list$clk                     = clk;
  assign free_list$free_call$000           = free_call$000;
  assign free_list$free_index$000          = free_index$000;
  assign free_list$release_mask            = dump_mux$mux_out;
  assign free_list$reset                   = reset;
  assign free_list$set_call                = set_call;
  assign free_list$set_state               = set_state;
  assign snapshot_packers$000$clk          = clk;
  assign snapshot_packers$000$pack_in_$000 = snapshots$000$dump_out$000;
  assign snapshot_packers$000$pack_in_$001 = snapshots$000$dump_out$001;
  assign snapshot_packers$000$reset        = reset;
  assign snapshot_packers$001$clk          = clk;
  assign snapshot_packers$001$pack_in_$000 = snapshots$001$dump_out$000;
  assign snapshot_packers$001$pack_in_$001 = snapshots$001$dump_out$001;
  assign snapshot_packers$001$reset        = reset;
  assign snapshots$000$clk                 = clk;
  assign snapshots$000$reset               = reset;
  assign snapshots$000$set_in_$000         = 1'd0;
  assign snapshots$000$set_in_$001         = 1'd0;
  assign snapshots$000$write_addr$000      = alloc_index$000;
  assign snapshots$000$write_call$000      = alloc_call$000;
  assign snapshots$000$write_data$000      = 1'd1;
  assign snapshots$001$clk                 = clk;
  assign snapshots$001$reset               = reset;
  assign snapshots$001$set_in_$000         = 1'd0;
  assign snapshots$001$set_in_$001         = 1'd0;
  assign snapshots$001$write_addr$000      = alloc_index$000;
  assign snapshots$001$write_call$000      = alloc_call$000;
  assign snapshots$001$write_data$000      = 1'd1;

  // array declarations
  logic    [   0:0] snapshots$set_call[0:1];
  assign snapshots$000$set_call = snapshots$set_call[  0];
  assign snapshots$001$set_call = snapshots$set_call[  1];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_reset_alloc_tracking_set_call(i=i):
  //         if s.reset_alloc_tracking_call and s.reset_alloc_tracking_target_id == i:
  //           s.snapshots[i].set_call.v = 1
  //         else:
  //           s.snapshots[i].set_call.v = 0

  // logic for handle_reset_alloc_tracking_set_call()
  always @ (*) begin
    if ((reset_alloc_tracking_call&&(reset_alloc_tracking_target_id == 0))) begin
      snapshots$set_call[0] = 1;
    end
    else begin
      snapshots$set_call[0] = 0;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_reset_alloc_tracking_set_call(i=i):
  //         if s.reset_alloc_tracking_call and s.reset_alloc_tracking_target_id == i:
  //           s.snapshots[i].set_call.v = 1
  //         else:
  //           s.snapshots[i].set_call.v = 0

  // logic for handle_reset_alloc_tracking_set_call()
  always @ (*) begin
    if ((reset_alloc_tracking_call&&(reset_alloc_tracking_target_id == 1))) begin
      snapshots$set_call[1] = 1;
    end
    else begin
      snapshots$set_call[1] = 0;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_revert_alloc():
  //       if s.reset_alloc_tracking_call and s.revert_allocs_call and s.reset_alloc_tracking_target_id == s.revert_allocs_source_id:
  //         s.free_list.release_call.v = 0
  //       else:
  //         s.free_list.release_call.v = s.revert_allocs_call

  // logic for handle_revert_alloc()
  always @ (*) begin
    if ((reset_alloc_tracking_call&&revert_allocs_call&&(reset_alloc_tracking_target_id == revert_allocs_source_id))) begin
      free_list$release_call = 0;
    end
    else begin
      free_list$release_call = revert_allocs_call;
    end
  end


endmodule // SnapshottingFreeList_0x64ee202bb6767a5b

//-----------------------------------------------------------------------------
// RegisterFile_0x6d9ba9c872129f4f
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.registerfile {"dtype": 1, "nregs": 2, "num_read_ports": 0, "num_write_ports": 1, "reset_values": null, "write_dump_bypass": true, "write_read_bypass": false}
// PyMTL: verilator_xinit = zeros
module RegisterFile_0x6d9ba9c872129f4f
(
  input  logic [   0:0] clk,
  output logic [   0:0] dump_out$000,
  output logic [   0:0] dump_out$001,
  input  logic [   0:0] reset,
  input  logic [   0:0] set_call,
  input  logic [   0:0] set_in_$000,
  input  logic [   0:0] set_in_$001,
  input  logic [   0:0] write_addr$000,
  input  logic [   0:0] write_call$000,
  input  logic [   0:0] write_data$000
);

  // logic declarations
  logic   [   0:0] write_inc$000;
  logic   [   0:0] write_inc$001;
  logic   [   0:0] after_set$000;
  logic   [   0:0] after_set$001;
  logic   [   0:0] regs$000;
  logic   [   0:0] regs$001;
  logic   [   0:0] after_write$000;
  logic   [   0:0] after_write$001;


  // signal connections
  assign dump_out$000 = after_write$000;
  assign dump_out$001 = after_write$001;

  // array declarations
  logic    [   0:0] after_set[0:1];
  assign after_set$000 = after_set[  0];
  assign after_set$001 = after_set[  1];
  logic    [   0:0] after_write[0:1];
  assign after_write$000 = after_write[  0];
  assign after_write$001 = after_write[  1];
  logic    [   0:0] regs[0:1];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  logic   [   0:0] set_in_[0:1];
  assign set_in_[  0] = set_in_$000;
  assign set_in_[  1] = set_in_$001;
  logic   [   0:0] write_addr[0:0];
  assign write_addr[  0] = write_addr$000;
  logic   [   0:0] write_call[0:0];
  assign write_call[  0] = write_call$000;
  logic   [   0:0] write_data[0:0];
  assign write_data[  0] = write_data$000;
  logic    [   0:0] write_inc[0:1];
  assign write_inc$000 = write_inc[  0];
  assign write_inc$001 = write_inc[  1];

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[0] <= 0;
    end
    else begin
      regs[0] <= after_set[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[1] <= 0;
    end
    else begin
      regs[1] <= after_set[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 0))) begin
      write_inc[0] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[0] = regs[0];
      end
      else begin
        write_inc[0] = write_inc[-2];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[0] = write_inc[0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[0] = set_in_[0];
    end
    else begin
      after_set[0] = after_write[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 1))) begin
      write_inc[1] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[1] = regs[1];
      end
      else begin
        write_inc[1] = write_inc[-1];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[1] = write_inc[1];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[1] = set_in_[1];
    end
    else begin
      after_set[1] = after_write[1];
    end
  end


endmodule // RegisterFile_0x6d9ba9c872129f4f

//-----------------------------------------------------------------------------
// Mux_0x7cc3cbcc1953dfea
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.mux {"dtype": 2, "nports": 2}
// PyMTL: verilator_xinit = zeros
module Mux_0x7cc3cbcc1953dfea
(
  input  logic [   0:0] clk,
  input  logic [   1:0] mux_in_$000,
  input  logic [   1:0] mux_in_$001,
  output logic  [   1:0] mux_out,
  input  logic [   0:0] mux_select,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nports = 2;


  // array declarations
  logic   [   1:0] mux_in_[0:1];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def select():
  //       assert s.mux_select < nports
  //       s.mux_out.v = s.mux_in_[s.mux_select]

  // logic for select()
  always @ (*) begin
    mux_out = mux_in_[mux_select];
  end


endmodule // Mux_0x7cc3cbcc1953dfea

//-----------------------------------------------------------------------------
// FreeList_0x260f6d53b9562731
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.freelist {"free_alloc_bypass": false, "nslots": 2, "num_alloc_ports": 1, "num_free_ports": 1, "release_alloc_bypass": false, "used_slots_initial": 0}
// PyMTL: verilator_xinit = zeros
module FreeList_0x260f6d53b9562731
(
  input  logic [   0:0] alloc_call$000,
  output logic [   0:0] alloc_index$000,
  output logic [   1:0] alloc_mask$000,
  output logic [   0:0] alloc_rdy$000,
  input  logic [   0:0] clk,
  input  logic [   0:0] free_call$000,
  input  logic [   0:0] free_index$000,
  input  logic [   0:0] release_call,
  input  logic [   1:0] release_mask,
  input  logic [   0:0] reset,
  input  logic [   0:0] set_call,
  input  logic [   1:0] set_state
);

  // logic declarations
  logic   [   1:0] free_masks$000;
  logic   [   1:0] free_masks$001;
  logic   [   1:0] alloc_inc$000;
  logic   [   1:0] alloc_inc$001;


  // register declarations
  logic    [   1:0] alloc_inc_base;
  logic    [   1:0] free_next;
  logic    [   1:0] free_next_base;
  logic    [   1:0] free_vector;

  // localparam declarations
  localparam num_alloc_ports = 1;
  localparam num_free_ports = 1;

  // free_encoders$000 temporaries
  logic   [   0:0] free_encoders$000$clk;
  logic   [   0:0] free_encoders$000$reset;
  logic   [   0:0] free_encoders$000$encode_number;
  logic   [   1:0] free_encoders$000$encode_onehot;

  OneHotEncoder_0x62af1c1ff9e32b51 free_encoders$000
  (
    .clk           ( free_encoders$000$clk ),
    .reset         ( free_encoders$000$reset ),
    .encode_number ( free_encoders$000$encode_number ),
    .encode_onehot ( free_encoders$000$encode_onehot )
  );

  // alloc_decoders$000 temporaries
  logic   [   0:0] alloc_decoders$000$clk;
  logic   [   0:0] alloc_decoders$000$reset;
  logic   [   1:0] alloc_decoders$000$decode_signal;
  logic   [   0:0] alloc_decoders$000$decode_valid;
  logic   [   0:0] alloc_decoders$000$decode_decoded;

  PriorityDecoder_0x86563bd99c43c59 alloc_decoders$000
  (
    .clk            ( alloc_decoders$000$clk ),
    .reset          ( alloc_decoders$000$reset ),
    .decode_signal  ( alloc_decoders$000$decode_signal ),
    .decode_valid   ( alloc_decoders$000$decode_valid ),
    .decode_decoded ( alloc_decoders$000$decode_decoded )
  );

  // alloc_encoders$000 temporaries
  logic   [   0:0] alloc_encoders$000$clk;
  logic   [   0:0] alloc_encoders$000$reset;
  logic   [   0:0] alloc_encoders$000$encode_number;
  logic   [   1:0] alloc_encoders$000$encode_onehot;

  OneHotEncoder_0x62af1c1ff9e32b51 alloc_encoders$000
  (
    .clk           ( alloc_encoders$000$clk ),
    .reset         ( alloc_encoders$000$reset ),
    .encode_number ( alloc_encoders$000$encode_number ),
    .encode_onehot ( alloc_encoders$000$encode_onehot )
  );

  // set_mux temporaries
  logic   [   1:0] set_mux$mux_in_$000;
  logic   [   1:0] set_mux$mux_in_$001;
  logic   [   0:0] set_mux$clk;
  logic   [   0:0] set_mux$reset;
  logic   [   0:0] set_mux$mux_select;
  logic   [   1:0] set_mux$mux_out;

  Mux_0x7cc3cbcc1953dfea set_mux
  (
    .mux_in_$000 ( set_mux$mux_in_$000 ),
    .mux_in_$001 ( set_mux$mux_in_$001 ),
    .clk         ( set_mux$clk ),
    .reset       ( set_mux$reset ),
    .mux_select  ( set_mux$mux_select ),
    .mux_out     ( set_mux$mux_out )
  );

  // signal connections
  assign alloc_decoders$000$clk           = clk;
  assign alloc_decoders$000$decode_signal = alloc_inc$000;
  assign alloc_decoders$000$reset         = reset;
  assign alloc_encoders$000$clk           = clk;
  assign alloc_encoders$000$encode_number = alloc_decoders$000$decode_decoded;
  assign alloc_encoders$000$reset         = reset;
  assign alloc_index$000                  = alloc_decoders$000$decode_decoded;
  assign alloc_mask$000                   = alloc_encoders$000$encode_onehot;
  assign alloc_rdy$000                    = alloc_decoders$000$decode_valid;
  assign free_encoders$000$clk            = clk;
  assign free_encoders$000$encode_number  = free_index$000;
  assign free_encoders$000$reset          = reset;
  assign free_masks$000                   = 2'd0;
  assign set_mux$clk                      = clk;
  assign set_mux$mux_in_$000              = free_next;
  assign set_mux$mux_in_$001              = set_state;
  assign set_mux$mux_select               = set_call;
  assign set_mux$reset                    = reset;

  // array declarations
  logic   [   0:0] alloc_call[0:0];
  assign alloc_call[  0] = alloc_call$000;
  logic   [   1:0] alloc_encoders$encode_onehot[0:0];
  assign alloc_encoders$encode_onehot[  0] = alloc_encoders$000$encode_onehot;
  logic    [   1:0] alloc_inc[0:1];
  assign alloc_inc$000 = alloc_inc[  0];
  assign alloc_inc$001 = alloc_inc[  1];
  logic   [   0:0] free_call[0:0];
  assign free_call[  0] = free_call$000;
  logic   [   1:0] free_encoders$encode_onehot[0:0];
  assign free_encoders$encode_onehot[  0] = free_encoders$000$encode_onehot;
  logic    [   1:0] free_masks[0:1];
  assign free_masks$000 = free_masks[  0];
  assign free_masks$001 = free_masks[  1];

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[0] <= 1;
    end
    else begin
      free_vector[0] <= set_mux$mux_out[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[1] <= 1;
    end
    else begin
      free_vector[1] <= set_mux$mux_out[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_free(n=i + 1, i=i):
  //         if s.free_call[i]:
  //           s.free_masks[n].v = s.free_masks[i] | s.free_encoders[i].encode_onehot
  //         else:
  //           s.free_masks[n].v = s.free_masks[i]

  // logic for handle_free()
  always @ (*) begin
    if (free_call[0]) begin
      free_masks[1] = (free_masks[0]|free_encoders$encode_onehot[0]);
    end
    else begin
      free_masks[1] = free_masks[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_alloc_inc_base():
  //         s.alloc_inc_base.v = s.free_vector

  // logic for compute_alloc_inc_base()
  always @ (*) begin
    alloc_inc_base = free_vector;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_alloc_inc_0():
  //         s.alloc_inc[0].v = s.alloc_inc_base

  // logic for compute_alloc_inc_0()
  always @ (*) begin
    alloc_inc[0] = alloc_inc_base;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_alloc(n=i + 1, i=i):
  //         if s.alloc_call[i]:
  //           s.alloc_inc[n].v = s.alloc_inc[i] & (
  //               ~s.alloc_encoders[i].encode_onehot)
  //         else:
  //           s.alloc_inc[n].v = s.alloc_inc[i]

  // logic for handle_alloc()
  always @ (*) begin
    if (alloc_call[0]) begin
      alloc_inc[1] = (alloc_inc[0]&~alloc_encoders$encode_onehot[0]);
    end
    else begin
      alloc_inc[1] = alloc_inc[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_free_next_base():
  //         if s.release_call:
  //           s.free_next_base.v = s.alloc_inc[num_alloc_ports] | s.release_mask
  //         else:
  //           s.free_next_base.v = s.alloc_inc[num_alloc_ports]

  // logic for compute_free_next_base()
  always @ (*) begin
    if (release_call) begin
      free_next_base = (alloc_inc[num_alloc_ports]|release_mask);
    end
    else begin
      free_next_base = alloc_inc[num_alloc_ports];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_free():
  //         s.free_next.v = s.free_next_base | s.free_masks[num_free_ports]

  // logic for compute_free()
  always @ (*) begin
    free_next = (free_next_base|free_masks[num_free_ports]);
  end


endmodule // FreeList_0x260f6d53b9562731

//-----------------------------------------------------------------------------
// AsynchronousRAM_0x49021b1555bbbcb6
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.async_ram {"interface": "read[2] (addr: Bits(6)) -> (data: Bits(1)); write[2] <C> (data: Bits(1), addr: Bits(6)) -> ()", "reset_values": 1}
// PyMTL: verilator_xinit = zeros
module AsynchronousRAM_0x49021b1555bbbcb6
(
  input  logic [   0:0] clk,
  input  logic [   5:0] read_addr$000,
  input  logic [   5:0] read_addr$001,
  output logic [   0:0] read_data$000,
  output logic [   0:0] read_data$001,
  input  logic [   0:0] reset,
  input  logic [   5:0] write_addr$000,
  input  logic [   5:0] write_addr$001,
  input  logic [   0:0] write_call$000,
  input  logic [   0:0] write_call$001,
  input  logic [   0:0] write_data$000,
  input  logic [   0:0] write_data$001
);

  // logic declarations
  logic   [   0:0] regs$000;
  logic   [   0:0] regs$001;
  logic   [   0:0] regs$002;
  logic   [   0:0] regs$003;
  logic   [   0:0] regs$004;
  logic   [   0:0] regs$005;
  logic   [   0:0] regs$006;
  logic   [   0:0] regs$007;
  logic   [   0:0] regs$008;
  logic   [   0:0] regs$009;
  logic   [   0:0] regs$010;
  logic   [   0:0] regs$011;
  logic   [   0:0] regs$012;
  logic   [   0:0] regs$013;
  logic   [   0:0] regs$014;
  logic   [   0:0] regs$015;
  logic   [   0:0] regs$016;
  logic   [   0:0] regs$017;
  logic   [   0:0] regs$018;
  logic   [   0:0] regs$019;
  logic   [   0:0] regs$020;
  logic   [   0:0] regs$021;
  logic   [   0:0] regs$022;
  logic   [   0:0] regs$023;
  logic   [   0:0] regs$024;
  logic   [   0:0] regs$025;
  logic   [   0:0] regs$026;
  logic   [   0:0] regs$027;
  logic   [   0:0] regs$028;
  logic   [   0:0] regs$029;
  logic   [   0:0] regs$030;
  logic   [   0:0] regs$031;
  logic   [   0:0] regs$032;
  logic   [   0:0] regs$033;
  logic   [   0:0] regs$034;
  logic   [   0:0] regs$035;
  logic   [   0:0] regs$036;
  logic   [   0:0] regs$037;
  logic   [   0:0] regs$038;
  logic   [   0:0] regs$039;
  logic   [   0:0] regs$040;
  logic   [   0:0] regs$041;
  logic   [   0:0] regs$042;
  logic   [   0:0] regs$043;
  logic   [   0:0] regs$044;
  logic   [   0:0] regs$045;
  logic   [   0:0] regs$046;
  logic   [   0:0] regs$047;
  logic   [   0:0] regs$048;
  logic   [   0:0] regs$049;
  logic   [   0:0] regs$050;
  logic   [   0:0] regs$051;
  logic   [   0:0] regs$052;
  logic   [   0:0] regs$053;
  logic   [   0:0] regs$054;
  logic   [   0:0] regs$055;
  logic   [   0:0] regs$056;
  logic   [   0:0] regs$057;
  logic   [   0:0] regs$058;
  logic   [   0:0] regs$059;
  logic   [   0:0] regs$060;
  logic   [   0:0] regs$061;
  logic   [   0:0] regs$062;
  logic   [   0:0] regs$063;


  // localparam declarations
  localparam num_read_ports = 2;
  localparam num_write_ports = 2;
  localparam nwords = 64;
  localparam reset_values = 1;

  // loop variable declarations
  integer i;


  // array declarations
  logic   [   5:0] read_addr[0:1];
  assign read_addr[  0] = read_addr$000;
  assign read_addr[  1] = read_addr$001;
  logic    [   0:0] read_data[0:1];
  assign read_data$000 = read_data[  0];
  assign read_data$001 = read_data[  1];
  logic    [   0:0] regs[0:63];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  assign regs$002 = regs[  2];
  assign regs$003 = regs[  3];
  assign regs$004 = regs[  4];
  assign regs$005 = regs[  5];
  assign regs$006 = regs[  6];
  assign regs$007 = regs[  7];
  assign regs$008 = regs[  8];
  assign regs$009 = regs[  9];
  assign regs$010 = regs[ 10];
  assign regs$011 = regs[ 11];
  assign regs$012 = regs[ 12];
  assign regs$013 = regs[ 13];
  assign regs$014 = regs[ 14];
  assign regs$015 = regs[ 15];
  assign regs$016 = regs[ 16];
  assign regs$017 = regs[ 17];
  assign regs$018 = regs[ 18];
  assign regs$019 = regs[ 19];
  assign regs$020 = regs[ 20];
  assign regs$021 = regs[ 21];
  assign regs$022 = regs[ 22];
  assign regs$023 = regs[ 23];
  assign regs$024 = regs[ 24];
  assign regs$025 = regs[ 25];
  assign regs$026 = regs[ 26];
  assign regs$027 = regs[ 27];
  assign regs$028 = regs[ 28];
  assign regs$029 = regs[ 29];
  assign regs$030 = regs[ 30];
  assign regs$031 = regs[ 31];
  assign regs$032 = regs[ 32];
  assign regs$033 = regs[ 33];
  assign regs$034 = regs[ 34];
  assign regs$035 = regs[ 35];
  assign regs$036 = regs[ 36];
  assign regs$037 = regs[ 37];
  assign regs$038 = regs[ 38];
  assign regs$039 = regs[ 39];
  assign regs$040 = regs[ 40];
  assign regs$041 = regs[ 41];
  assign regs$042 = regs[ 42];
  assign regs$043 = regs[ 43];
  assign regs$044 = regs[ 44];
  assign regs$045 = regs[ 45];
  assign regs$046 = regs[ 46];
  assign regs$047 = regs[ 47];
  assign regs$048 = regs[ 48];
  assign regs$049 = regs[ 49];
  assign regs$050 = regs[ 50];
  assign regs$051 = regs[ 51];
  assign regs$052 = regs[ 52];
  assign regs$053 = regs[ 53];
  assign regs$054 = regs[ 54];
  assign regs$055 = regs[ 55];
  assign regs$056 = regs[ 56];
  assign regs$057 = regs[ 57];
  assign regs$058 = regs[ 58];
  assign regs$059 = regs[ 59];
  assign regs$060 = regs[ 60];
  assign regs$061 = regs[ 61];
  assign regs$062 = regs[ 62];
  assign regs$063 = regs[ 63];
  logic   [   5:0] write_addr[0:1];
  assign write_addr[  0] = write_addr$000;
  assign write_addr[  1] = write_addr$001;
  logic   [   0:0] write_call[0:1];
  assign write_call[  0] = write_call$000;
  assign write_call[  1] = write_call$001;
  logic   [   0:0] write_data[0:1];
  assign write_data[  0] = write_data$000;
  assign write_data[  1] = write_data$001;

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def handle_writes():
  //         if s.reset:
  //           for i in range(nwords):
  //             s.regs[i].n = reset_values
  //         else:
  //           for i in range(num_write_ports):
  //             if s.write_call[i]:
  //               s.regs[s.write_addr[i]].n = s.write_data[i]

  // logic for handle_writes()
  always @ (posedge clk) begin
    if (reset) begin
      for (i=0; i < nwords; i=i+1)
      begin
        regs[i] <= reset_values;
      end
    end
    else begin
      for (i=0; i < num_write_ports; i=i+1)
      begin
        if (write_call[i]) begin
          regs[write_addr[i]] <= write_data[i];
        end
        else begin
        end
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_reads():
  //         for i in range(num_read_ports):
  //           s.read_data[i].v = s.regs[s.read_addr[i]]

  // logic for handle_reads()
  always @ (*) begin
    for (i=0; i < num_read_ports; i=i+1)
    begin
      read_data[i] = regs[read_addr[i]];
    end
  end


endmodule // AsynchronousRAM_0x49021b1555bbbcb6

//-----------------------------------------------------------------------------
// Mux_0x183cf582fc8d227d
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.mux {"dtype": 1, "nports": 2}
// PyMTL: verilator_xinit = zeros
module Mux_0x183cf582fc8d227d
(
  input  logic [   0:0] clk,
  input  logic [   0:0] mux_in_$000,
  input  logic [   0:0] mux_in_$001,
  output logic  [   0:0] mux_out,
  input  logic [   0:0] mux_select,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nports = 2;


  // array declarations
  logic   [   0:0] mux_in_[0:1];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def select():
  //       assert s.mux_select < nports
  //       s.mux_out.v = s.mux_in_[s.mux_select]

  // logic for select()
  always @ (*) begin
    mux_out = mux_in_[mux_select];
  end


endmodule // Mux_0x183cf582fc8d227d

//-----------------------------------------------------------------------------
// Packer_0x5417ceb8bd59f204
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.packers {"dtype": 1, "nports": 63}
// PyMTL: verilator_xinit = zeros
module Packer_0x5417ceb8bd59f204
(
  input  logic [   0:0] clk,
  input  logic [   0:0] pack_in_$000,
  input  logic [   0:0] pack_in_$010,
  input  logic [   0:0] pack_in_$011,
  input  logic [   0:0] pack_in_$012,
  input  logic [   0:0] pack_in_$013,
  input  logic [   0:0] pack_in_$014,
  input  logic [   0:0] pack_in_$015,
  input  logic [   0:0] pack_in_$016,
  input  logic [   0:0] pack_in_$017,
  input  logic [   0:0] pack_in_$018,
  input  logic [   0:0] pack_in_$019,
  input  logic [   0:0] pack_in_$001,
  input  logic [   0:0] pack_in_$020,
  input  logic [   0:0] pack_in_$021,
  input  logic [   0:0] pack_in_$022,
  input  logic [   0:0] pack_in_$023,
  input  logic [   0:0] pack_in_$024,
  input  logic [   0:0] pack_in_$025,
  input  logic [   0:0] pack_in_$026,
  input  logic [   0:0] pack_in_$027,
  input  logic [   0:0] pack_in_$028,
  input  logic [   0:0] pack_in_$029,
  input  logic [   0:0] pack_in_$002,
  input  logic [   0:0] pack_in_$030,
  input  logic [   0:0] pack_in_$031,
  input  logic [   0:0] pack_in_$032,
  input  logic [   0:0] pack_in_$033,
  input  logic [   0:0] pack_in_$034,
  input  logic [   0:0] pack_in_$035,
  input  logic [   0:0] pack_in_$036,
  input  logic [   0:0] pack_in_$037,
  input  logic [   0:0] pack_in_$038,
  input  logic [   0:0] pack_in_$039,
  input  logic [   0:0] pack_in_$003,
  input  logic [   0:0] pack_in_$040,
  input  logic [   0:0] pack_in_$041,
  input  logic [   0:0] pack_in_$042,
  input  logic [   0:0] pack_in_$043,
  input  logic [   0:0] pack_in_$044,
  input  logic [   0:0] pack_in_$045,
  input  logic [   0:0] pack_in_$046,
  input  logic [   0:0] pack_in_$047,
  input  logic [   0:0] pack_in_$048,
  input  logic [   0:0] pack_in_$049,
  input  logic [   0:0] pack_in_$004,
  input  logic [   0:0] pack_in_$050,
  input  logic [   0:0] pack_in_$051,
  input  logic [   0:0] pack_in_$052,
  input  logic [   0:0] pack_in_$053,
  input  logic [   0:0] pack_in_$054,
  input  logic [   0:0] pack_in_$055,
  input  logic [   0:0] pack_in_$056,
  input  logic [   0:0] pack_in_$057,
  input  logic [   0:0] pack_in_$058,
  input  logic [   0:0] pack_in_$059,
  input  logic [   0:0] pack_in_$005,
  input  logic [   0:0] pack_in_$060,
  input  logic [   0:0] pack_in_$061,
  input  logic [   0:0] pack_in_$062,
  input  logic [   0:0] pack_in_$006,
  input  logic [   0:0] pack_in_$007,
  input  logic [   0:0] pack_in_$008,
  input  logic [   0:0] pack_in_$009,
  output logic  [  62:0] pack_packed,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nbits = 1;


  // array declarations
  logic   [   0:0] pack_in_[0:62];
  assign pack_in_[  0] = pack_in_$000;
  assign pack_in_[  1] = pack_in_$001;
  assign pack_in_[  2] = pack_in_$002;
  assign pack_in_[  3] = pack_in_$003;
  assign pack_in_[  4] = pack_in_$004;
  assign pack_in_[  5] = pack_in_$005;
  assign pack_in_[  6] = pack_in_$006;
  assign pack_in_[  7] = pack_in_$007;
  assign pack_in_[  8] = pack_in_$008;
  assign pack_in_[  9] = pack_in_$009;
  assign pack_in_[ 10] = pack_in_$010;
  assign pack_in_[ 11] = pack_in_$011;
  assign pack_in_[ 12] = pack_in_$012;
  assign pack_in_[ 13] = pack_in_$013;
  assign pack_in_[ 14] = pack_in_$014;
  assign pack_in_[ 15] = pack_in_$015;
  assign pack_in_[ 16] = pack_in_$016;
  assign pack_in_[ 17] = pack_in_$017;
  assign pack_in_[ 18] = pack_in_$018;
  assign pack_in_[ 19] = pack_in_$019;
  assign pack_in_[ 20] = pack_in_$020;
  assign pack_in_[ 21] = pack_in_$021;
  assign pack_in_[ 22] = pack_in_$022;
  assign pack_in_[ 23] = pack_in_$023;
  assign pack_in_[ 24] = pack_in_$024;
  assign pack_in_[ 25] = pack_in_$025;
  assign pack_in_[ 26] = pack_in_$026;
  assign pack_in_[ 27] = pack_in_$027;
  assign pack_in_[ 28] = pack_in_$028;
  assign pack_in_[ 29] = pack_in_$029;
  assign pack_in_[ 30] = pack_in_$030;
  assign pack_in_[ 31] = pack_in_$031;
  assign pack_in_[ 32] = pack_in_$032;
  assign pack_in_[ 33] = pack_in_$033;
  assign pack_in_[ 34] = pack_in_$034;
  assign pack_in_[ 35] = pack_in_$035;
  assign pack_in_[ 36] = pack_in_$036;
  assign pack_in_[ 37] = pack_in_$037;
  assign pack_in_[ 38] = pack_in_$038;
  assign pack_in_[ 39] = pack_in_$039;
  assign pack_in_[ 40] = pack_in_$040;
  assign pack_in_[ 41] = pack_in_$041;
  assign pack_in_[ 42] = pack_in_$042;
  assign pack_in_[ 43] = pack_in_$043;
  assign pack_in_[ 44] = pack_in_$044;
  assign pack_in_[ 45] = pack_in_$045;
  assign pack_in_[ 46] = pack_in_$046;
  assign pack_in_[ 47] = pack_in_$047;
  assign pack_in_[ 48] = pack_in_$048;
  assign pack_in_[ 49] = pack_in_$049;
  assign pack_in_[ 50] = pack_in_$050;
  assign pack_in_[ 51] = pack_in_$051;
  assign pack_in_[ 52] = pack_in_$052;
  assign pack_in_[ 53] = pack_in_$053;
  assign pack_in_[ 54] = pack_in_$054;
  assign pack_in_[ 55] = pack_in_$055;
  assign pack_in_[ 56] = pack_in_$056;
  assign pack_in_[ 57] = pack_in_$057;
  assign pack_in_[ 58] = pack_in_$058;
  assign pack_in_[ 59] = pack_in_$059;
  assign pack_in_[ 60] = pack_in_$060;
  assign pack_in_[ 61] = pack_in_$061;
  assign pack_in_[ 62] = pack_in_$062;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(1)-1:0] = pack_in_[0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(2)-1:1] = pack_in_[1];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(3)-1:2] = pack_in_[2];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(4)-1:3] = pack_in_[3];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(5)-1:4] = pack_in_[4];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(6)-1:5] = pack_in_[5];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(7)-1:6] = pack_in_[6];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(8)-1:7] = pack_in_[7];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(9)-1:8] = pack_in_[8];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(10)-1:9] = pack_in_[9];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(11)-1:10] = pack_in_[10];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(12)-1:11] = pack_in_[11];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(13)-1:12] = pack_in_[12];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(14)-1:13] = pack_in_[13];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(15)-1:14] = pack_in_[14];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(16)-1:15] = pack_in_[15];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(17)-1:16] = pack_in_[16];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(18)-1:17] = pack_in_[17];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(19)-1:18] = pack_in_[18];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(20)-1:19] = pack_in_[19];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(21)-1:20] = pack_in_[20];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(22)-1:21] = pack_in_[21];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(23)-1:22] = pack_in_[22];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(24)-1:23] = pack_in_[23];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(25)-1:24] = pack_in_[24];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(26)-1:25] = pack_in_[25];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(27)-1:26] = pack_in_[26];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(28)-1:27] = pack_in_[27];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(29)-1:28] = pack_in_[28];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(30)-1:29] = pack_in_[29];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(31)-1:30] = pack_in_[30];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(32)-1:31] = pack_in_[31];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(33)-1:32] = pack_in_[32];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(34)-1:33] = pack_in_[33];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(35)-1:34] = pack_in_[34];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(36)-1:35] = pack_in_[35];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(37)-1:36] = pack_in_[36];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(38)-1:37] = pack_in_[37];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(39)-1:38] = pack_in_[38];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(40)-1:39] = pack_in_[39];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(41)-1:40] = pack_in_[40];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(42)-1:41] = pack_in_[41];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(43)-1:42] = pack_in_[42];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(44)-1:43] = pack_in_[43];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(45)-1:44] = pack_in_[44];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(46)-1:45] = pack_in_[45];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(47)-1:46] = pack_in_[46];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(48)-1:47] = pack_in_[47];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(49)-1:48] = pack_in_[48];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(50)-1:49] = pack_in_[49];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(51)-1:50] = pack_in_[50];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(52)-1:51] = pack_in_[51];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(53)-1:52] = pack_in_[52];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(54)-1:53] = pack_in_[53];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(55)-1:54] = pack_in_[54];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(56)-1:55] = pack_in_[55];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(57)-1:56] = pack_in_[56];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(58)-1:57] = pack_in_[57];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(59)-1:58] = pack_in_[58];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(60)-1:59] = pack_in_[59];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(61)-1:60] = pack_in_[60];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(62)-1:61] = pack_in_[61];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pack(i=i,
  //                start=i * s.interface.Data.nbits,
  //                end=(i + 1) * s.interface.Data.nbits):
  //         s.pack_packed[start:end].v = s.pack_in_[i]

  // logic for pack()
  always @ (*) begin
    pack_packed[(63)-1:62] = pack_in_[62];
  end


endmodule // Packer_0x5417ceb8bd59f204

//-----------------------------------------------------------------------------
// RenameTable_0x2b84c99320ad3cb1
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.renametable {"const_zero": true, "initial_map": [0, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30], "naregs": 32, "npregs": 64, "nsnapshots": 2, "num_lookup_ports": 2, "num_update_ports": 1}
// PyMTL: verilator_xinit = zeros
module RenameTable_0x2b84c99320ad3cb1
(
  input  logic [   0:0] clk,
  input  logic [   4:0] lookup_areg$000,
  input  logic [   4:0] lookup_areg$001,
  output logic [   5:0] lookup_preg$000,
  output logic [   5:0] lookup_preg$001,
  input  logic [   0:0] reset,
  input  logic [   0:0] restore_call,
  input  logic [   0:0] restore_source_id,
  input  logic [   0:0] set_call,
  input  logic [   5:0] set_in_$000,
  input  logic [   5:0] set_in_$010,
  input  logic [   5:0] set_in_$011,
  input  logic [   5:0] set_in_$012,
  input  logic [   5:0] set_in_$013,
  input  logic [   5:0] set_in_$014,
  input  logic [   5:0] set_in_$015,
  input  logic [   5:0] set_in_$016,
  input  logic [   5:0] set_in_$017,
  input  logic [   5:0] set_in_$018,
  input  logic [   5:0] set_in_$019,
  input  logic [   5:0] set_in_$001,
  input  logic [   5:0] set_in_$020,
  input  logic [   5:0] set_in_$021,
  input  logic [   5:0] set_in_$022,
  input  logic [   5:0] set_in_$023,
  input  logic [   5:0] set_in_$024,
  input  logic [   5:0] set_in_$025,
  input  logic [   5:0] set_in_$026,
  input  logic [   5:0] set_in_$027,
  input  logic [   5:0] set_in_$028,
  input  logic [   5:0] set_in_$029,
  input  logic [   5:0] set_in_$002,
  input  logic [   5:0] set_in_$030,
  input  logic [   5:0] set_in_$031,
  input  logic [   5:0] set_in_$003,
  input  logic [   5:0] set_in_$004,
  input  logic [   5:0] set_in_$005,
  input  logic [   5:0] set_in_$006,
  input  logic [   5:0] set_in_$007,
  input  logic [   5:0] set_in_$008,
  input  logic [   5:0] set_in_$009,
  input  logic [   0:0] snapshot_call,
  input  logic [   0:0] snapshot_target_id,
  input  logic [   4:0] update_areg$000,
  input  logic [   0:0] update_call$000,
  input  logic [   5:0] update_preg$000
);

  // localparam declarations
  localparam ZERO_TAG = 6'd63;

  // rename_table temporaries
  logic   [   0:0] rename_table$snapshot_call;
  logic   [   5:0] rename_table$set_in_$000;
  logic   [   5:0] rename_table$set_in_$001;
  logic   [   5:0] rename_table$set_in_$002;
  logic   [   5:0] rename_table$set_in_$003;
  logic   [   5:0] rename_table$set_in_$004;
  logic   [   5:0] rename_table$set_in_$005;
  logic   [   5:0] rename_table$set_in_$006;
  logic   [   5:0] rename_table$set_in_$007;
  logic   [   5:0] rename_table$set_in_$008;
  logic   [   5:0] rename_table$set_in_$009;
  logic   [   5:0] rename_table$set_in_$010;
  logic   [   5:0] rename_table$set_in_$011;
  logic   [   5:0] rename_table$set_in_$012;
  logic   [   5:0] rename_table$set_in_$013;
  logic   [   5:0] rename_table$set_in_$014;
  logic   [   5:0] rename_table$set_in_$015;
  logic   [   5:0] rename_table$set_in_$016;
  logic   [   5:0] rename_table$set_in_$017;
  logic   [   5:0] rename_table$set_in_$018;
  logic   [   5:0] rename_table$set_in_$019;
  logic   [   5:0] rename_table$set_in_$020;
  logic   [   5:0] rename_table$set_in_$021;
  logic   [   5:0] rename_table$set_in_$022;
  logic   [   5:0] rename_table$set_in_$023;
  logic   [   5:0] rename_table$set_in_$024;
  logic   [   5:0] rename_table$set_in_$025;
  logic   [   5:0] rename_table$set_in_$026;
  logic   [   5:0] rename_table$set_in_$027;
  logic   [   5:0] rename_table$set_in_$028;
  logic   [   5:0] rename_table$set_in_$029;
  logic   [   5:0] rename_table$set_in_$030;
  logic   [   5:0] rename_table$set_in_$031;
  logic   [   0:0] rename_table$set_call;
  logic   [   0:0] rename_table$restore_source_id;
  logic   [   0:0] rename_table$restore_call;
  logic   [   0:0] rename_table$clk;
  logic   [   4:0] rename_table$write_addr$000;
  logic   [   4:0] rename_table$read_addr$000;
  logic   [   4:0] rename_table$read_addr$001;
  logic   [   0:0] rename_table$write_call$000;
  logic   [   0:0] rename_table$snapshot_target_id;
  logic   [   5:0] rename_table$write_data$000;
  logic   [   0:0] rename_table$reset;
  logic   [   5:0] rename_table$read_data$000;
  logic   [   5:0] rename_table$read_data$001;

  SnapshottingRegisterFile_0x66bdadc3daaa062 rename_table
  (
    .snapshot_call      ( rename_table$snapshot_call ),
    .set_in_$000        ( rename_table$set_in_$000 ),
    .set_in_$001        ( rename_table$set_in_$001 ),
    .set_in_$002        ( rename_table$set_in_$002 ),
    .set_in_$003        ( rename_table$set_in_$003 ),
    .set_in_$004        ( rename_table$set_in_$004 ),
    .set_in_$005        ( rename_table$set_in_$005 ),
    .set_in_$006        ( rename_table$set_in_$006 ),
    .set_in_$007        ( rename_table$set_in_$007 ),
    .set_in_$008        ( rename_table$set_in_$008 ),
    .set_in_$009        ( rename_table$set_in_$009 ),
    .set_in_$010        ( rename_table$set_in_$010 ),
    .set_in_$011        ( rename_table$set_in_$011 ),
    .set_in_$012        ( rename_table$set_in_$012 ),
    .set_in_$013        ( rename_table$set_in_$013 ),
    .set_in_$014        ( rename_table$set_in_$014 ),
    .set_in_$015        ( rename_table$set_in_$015 ),
    .set_in_$016        ( rename_table$set_in_$016 ),
    .set_in_$017        ( rename_table$set_in_$017 ),
    .set_in_$018        ( rename_table$set_in_$018 ),
    .set_in_$019        ( rename_table$set_in_$019 ),
    .set_in_$020        ( rename_table$set_in_$020 ),
    .set_in_$021        ( rename_table$set_in_$021 ),
    .set_in_$022        ( rename_table$set_in_$022 ),
    .set_in_$023        ( rename_table$set_in_$023 ),
    .set_in_$024        ( rename_table$set_in_$024 ),
    .set_in_$025        ( rename_table$set_in_$025 ),
    .set_in_$026        ( rename_table$set_in_$026 ),
    .set_in_$027        ( rename_table$set_in_$027 ),
    .set_in_$028        ( rename_table$set_in_$028 ),
    .set_in_$029        ( rename_table$set_in_$029 ),
    .set_in_$030        ( rename_table$set_in_$030 ),
    .set_in_$031        ( rename_table$set_in_$031 ),
    .set_call           ( rename_table$set_call ),
    .restore_source_id  ( rename_table$restore_source_id ),
    .restore_call       ( rename_table$restore_call ),
    .clk                ( rename_table$clk ),
    .write_addr$000     ( rename_table$write_addr$000 ),
    .read_addr$000      ( rename_table$read_addr$000 ),
    .read_addr$001      ( rename_table$read_addr$001 ),
    .write_call$000     ( rename_table$write_call$000 ),
    .snapshot_target_id ( rename_table$snapshot_target_id ),
    .write_data$000     ( rename_table$write_data$000 ),
    .reset              ( rename_table$reset ),
    .read_data$000      ( rename_table$read_data$000 ),
    .read_data$001      ( rename_table$read_data$001 )
  );

  // signal connections
  assign rename_table$clk                = clk;
  assign rename_table$read_addr$000      = lookup_areg$000;
  assign rename_table$read_addr$001      = lookup_areg$001;
  assign rename_table$reset              = reset;
  assign rename_table$restore_call       = restore_call;
  assign rename_table$restore_source_id  = restore_source_id;
  assign rename_table$set_call           = set_call;
  assign rename_table$set_in_$000        = set_in_$000;
  assign rename_table$set_in_$001        = set_in_$001;
  assign rename_table$set_in_$002        = set_in_$002;
  assign rename_table$set_in_$003        = set_in_$003;
  assign rename_table$set_in_$004        = set_in_$004;
  assign rename_table$set_in_$005        = set_in_$005;
  assign rename_table$set_in_$006        = set_in_$006;
  assign rename_table$set_in_$007        = set_in_$007;
  assign rename_table$set_in_$008        = set_in_$008;
  assign rename_table$set_in_$009        = set_in_$009;
  assign rename_table$set_in_$010        = set_in_$010;
  assign rename_table$set_in_$011        = set_in_$011;
  assign rename_table$set_in_$012        = set_in_$012;
  assign rename_table$set_in_$013        = set_in_$013;
  assign rename_table$set_in_$014        = set_in_$014;
  assign rename_table$set_in_$015        = set_in_$015;
  assign rename_table$set_in_$016        = set_in_$016;
  assign rename_table$set_in_$017        = set_in_$017;
  assign rename_table$set_in_$018        = set_in_$018;
  assign rename_table$set_in_$019        = set_in_$019;
  assign rename_table$set_in_$020        = set_in_$020;
  assign rename_table$set_in_$021        = set_in_$021;
  assign rename_table$set_in_$022        = set_in_$022;
  assign rename_table$set_in_$023        = set_in_$023;
  assign rename_table$set_in_$024        = set_in_$024;
  assign rename_table$set_in_$025        = set_in_$025;
  assign rename_table$set_in_$026        = set_in_$026;
  assign rename_table$set_in_$027        = set_in_$027;
  assign rename_table$set_in_$028        = set_in_$028;
  assign rename_table$set_in_$029        = set_in_$029;
  assign rename_table$set_in_$030        = set_in_$030;
  assign rename_table$set_in_$031        = set_in_$031;
  assign rename_table$snapshot_call      = snapshot_call;
  assign rename_table$snapshot_target_id = snapshot_target_id;
  assign rename_table$write_addr$000     = update_areg$000;
  assign rename_table$write_data$000     = update_preg$000;

  // array declarations
  logic   [   4:0] lookup_areg[0:1];
  assign lookup_areg[  0] = lookup_areg$000;
  assign lookup_areg[  1] = lookup_areg$001;
  logic    [   5:0] lookup_preg[0:1];
  assign lookup_preg$000 = lookup_preg[  0];
  assign lookup_preg$001 = lookup_preg[  1];
  logic   [   5:0] rename_table$read_data[0:1];
  assign rename_table$read_data[  0] = rename_table$read_data$000;
  assign rename_table$read_data[  1] = rename_table$read_data$001;
  logic    [   0:0] rename_table$write_call[0:0];
  assign rename_table$write_call$000 = rename_table$write_call[  0];
  logic   [   4:0] update_areg[0:0];
  assign update_areg[  0] = update_areg$000;
  logic   [   0:0] update_call[0:0];
  assign update_call[  0] = update_call$000;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_zero_read(i=i):
  //           if s.lookup_areg[i] == 0:
  //             s.lookup_preg[i].v = s.ZERO_TAG
  //           else:
  //             s.lookup_preg[i].v = s.rename_table.read_data[i]

  // logic for handle_zero_read()
  always @ (*) begin
    if ((lookup_areg[0] == 0)) begin
      lookup_preg[0] = ZERO_TAG;
    end
    else begin
      lookup_preg[0] = rename_table$read_data[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_zero_read(i=i):
  //           if s.lookup_areg[i] == 0:
  //             s.lookup_preg[i].v = s.ZERO_TAG
  //           else:
  //             s.lookup_preg[i].v = s.rename_table.read_data[i]

  // logic for handle_zero_read()
  always @ (*) begin
    if ((lookup_areg[1] == 0)) begin
      lookup_preg[1] = ZERO_TAG;
    end
    else begin
      lookup_preg[1] = rename_table$read_data[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_zero_write(i=i):
  //           if s.update_areg[i] == 0:
  //             s.rename_table.write_call[i].v = 0
  //           else:
  //             s.rename_table.write_call[i].v = s.update_call[i]

  // logic for handle_zero_write()
  always @ (*) begin
    if ((update_areg[0] == 0)) begin
      rename_table$write_call[0] = 0;
    end
    else begin
      rename_table$write_call[0] = update_call[0];
    end
  end


endmodule // RenameTable_0x2b84c99320ad3cb1

//-----------------------------------------------------------------------------
// SnapshottingRegisterFile_0x66bdadc3daaa062
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.snapshotting_registerfile {"dtype": 6, "nregs": 32, "nsnapshots": 2, "num_read_ports": 2, "num_write_ports": 1, "reset_values": [0, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30], "write_read_bypass": false, "write_snapshot_bypass": true}
// PyMTL: verilator_xinit = zeros
module SnapshottingRegisterFile_0x66bdadc3daaa062
(
  input  logic [   0:0] clk,
  input  logic [   4:0] read_addr$000,
  input  logic [   4:0] read_addr$001,
  output logic [   5:0] read_data$000,
  output logic [   5:0] read_data$001,
  input  logic [   0:0] reset,
  input  logic [   0:0] restore_call,
  input  logic [   0:0] restore_source_id,
  input  logic [   0:0] set_call,
  input  logic [   5:0] set_in_$000,
  input  logic [   5:0] set_in_$010,
  input  logic [   5:0] set_in_$011,
  input  logic [   5:0] set_in_$012,
  input  logic [   5:0] set_in_$013,
  input  logic [   5:0] set_in_$014,
  input  logic [   5:0] set_in_$015,
  input  logic [   5:0] set_in_$016,
  input  logic [   5:0] set_in_$017,
  input  logic [   5:0] set_in_$018,
  input  logic [   5:0] set_in_$019,
  input  logic [   5:0] set_in_$001,
  input  logic [   5:0] set_in_$020,
  input  logic [   5:0] set_in_$021,
  input  logic [   5:0] set_in_$022,
  input  logic [   5:0] set_in_$023,
  input  logic [   5:0] set_in_$024,
  input  logic [   5:0] set_in_$025,
  input  logic [   5:0] set_in_$026,
  input  logic [   5:0] set_in_$027,
  input  logic [   5:0] set_in_$028,
  input  logic [   5:0] set_in_$029,
  input  logic [   5:0] set_in_$002,
  input  logic [   5:0] set_in_$030,
  input  logic [   5:0] set_in_$031,
  input  logic [   5:0] set_in_$003,
  input  logic [   5:0] set_in_$004,
  input  logic [   5:0] set_in_$005,
  input  logic [   5:0] set_in_$006,
  input  logic [   5:0] set_in_$007,
  input  logic [   5:0] set_in_$008,
  input  logic [   5:0] set_in_$009,
  input  logic [   0:0] snapshot_call,
  input  logic [   0:0] snapshot_target_id,
  input  logic [   4:0] write_addr$000,
  input  logic [   0:0] write_call$000,
  input  logic [   5:0] write_data$000
);

  // logic declarations
  logic   [   5:0] restore_vector$000;
  logic   [   5:0] restore_vector$001;
  logic   [   5:0] restore_vector$002;
  logic   [   5:0] restore_vector$003;
  logic   [   5:0] restore_vector$004;
  logic   [   5:0] restore_vector$005;
  logic   [   5:0] restore_vector$006;
  logic   [   5:0] restore_vector$007;
  logic   [   5:0] restore_vector$008;
  logic   [   5:0] restore_vector$009;
  logic   [   5:0] restore_vector$010;
  logic   [   5:0] restore_vector$011;
  logic   [   5:0] restore_vector$012;
  logic   [   5:0] restore_vector$013;
  logic   [   5:0] restore_vector$014;
  logic   [   5:0] restore_vector$015;
  logic   [   5:0] restore_vector$016;
  logic   [   5:0] restore_vector$017;
  logic   [   5:0] restore_vector$018;
  logic   [   5:0] restore_vector$019;
  logic   [   5:0] restore_vector$020;
  logic   [   5:0] restore_vector$021;
  logic   [   5:0] restore_vector$022;
  logic   [   5:0] restore_vector$023;
  logic   [   5:0] restore_vector$024;
  logic   [   5:0] restore_vector$025;
  logic   [   5:0] restore_vector$026;
  logic   [   5:0] restore_vector$027;
  logic   [   5:0] restore_vector$028;
  logic   [   5:0] restore_vector$029;
  logic   [   5:0] restore_vector$030;
  logic   [   5:0] restore_vector$031;
  logic   [   5:0] set_vector$000;
  logic   [   5:0] set_vector$001;
  logic   [   5:0] set_vector$002;
  logic   [   5:0] set_vector$003;
  logic   [   5:0] set_vector$004;
  logic   [   5:0] set_vector$005;
  logic   [   5:0] set_vector$006;
  logic   [   5:0] set_vector$007;
  logic   [   5:0] set_vector$008;
  logic   [   5:0] set_vector$009;
  logic   [   5:0] set_vector$010;
  logic   [   5:0] set_vector$011;
  logic   [   5:0] set_vector$012;
  logic   [   5:0] set_vector$013;
  logic   [   5:0] set_vector$014;
  logic   [   5:0] set_vector$015;
  logic   [   5:0] set_vector$016;
  logic   [   5:0] set_vector$017;
  logic   [   5:0] set_vector$018;
  logic   [   5:0] set_vector$019;
  logic   [   5:0] set_vector$020;
  logic   [   5:0] set_vector$021;
  logic   [   5:0] set_vector$022;
  logic   [   5:0] set_vector$023;
  logic   [   5:0] set_vector$024;
  logic   [   5:0] set_vector$025;
  logic   [   5:0] set_vector$026;
  logic   [   5:0] set_vector$027;
  logic   [   5:0] set_vector$028;
  logic   [   5:0] set_vector$029;
  logic   [   5:0] set_vector$030;
  logic   [   5:0] set_vector$031;


  // register declarations
  logic    [   0:0] should_restore;
  logic    [   0:0] should_set;

  // regs temporaries
  logic   [   5:0] regs$set_in_$000;
  logic   [   5:0] regs$set_in_$001;
  logic   [   5:0] regs$set_in_$002;
  logic   [   5:0] regs$set_in_$003;
  logic   [   5:0] regs$set_in_$004;
  logic   [   5:0] regs$set_in_$005;
  logic   [   5:0] regs$set_in_$006;
  logic   [   5:0] regs$set_in_$007;
  logic   [   5:0] regs$set_in_$008;
  logic   [   5:0] regs$set_in_$009;
  logic   [   5:0] regs$set_in_$010;
  logic   [   5:0] regs$set_in_$011;
  logic   [   5:0] regs$set_in_$012;
  logic   [   5:0] regs$set_in_$013;
  logic   [   5:0] regs$set_in_$014;
  logic   [   5:0] regs$set_in_$015;
  logic   [   5:0] regs$set_in_$016;
  logic   [   5:0] regs$set_in_$017;
  logic   [   5:0] regs$set_in_$018;
  logic   [   5:0] regs$set_in_$019;
  logic   [   5:0] regs$set_in_$020;
  logic   [   5:0] regs$set_in_$021;
  logic   [   5:0] regs$set_in_$022;
  logic   [   5:0] regs$set_in_$023;
  logic   [   5:0] regs$set_in_$024;
  logic   [   5:0] regs$set_in_$025;
  logic   [   5:0] regs$set_in_$026;
  logic   [   5:0] regs$set_in_$027;
  logic   [   5:0] regs$set_in_$028;
  logic   [   5:0] regs$set_in_$029;
  logic   [   5:0] regs$set_in_$030;
  logic   [   5:0] regs$set_in_$031;
  logic   [   0:0] regs$set_call;
  logic   [   0:0] regs$clk;
  logic   [   4:0] regs$write_addr$000;
  logic   [   4:0] regs$read_addr$000;
  logic   [   4:0] regs$read_addr$001;
  logic   [   0:0] regs$write_call$000;
  logic   [   5:0] regs$write_data$000;
  logic   [   0:0] regs$reset;
  logic   [   5:0] regs$read_data$000;
  logic   [   5:0] regs$read_data$001;
  logic   [   5:0] regs$dump_out$000;
  logic   [   5:0] regs$dump_out$001;
  logic   [   5:0] regs$dump_out$002;
  logic   [   5:0] regs$dump_out$003;
  logic   [   5:0] regs$dump_out$004;
  logic   [   5:0] regs$dump_out$005;
  logic   [   5:0] regs$dump_out$006;
  logic   [   5:0] regs$dump_out$007;
  logic   [   5:0] regs$dump_out$008;
  logic   [   5:0] regs$dump_out$009;
  logic   [   5:0] regs$dump_out$010;
  logic   [   5:0] regs$dump_out$011;
  logic   [   5:0] regs$dump_out$012;
  logic   [   5:0] regs$dump_out$013;
  logic   [   5:0] regs$dump_out$014;
  logic   [   5:0] regs$dump_out$015;
  logic   [   5:0] regs$dump_out$016;
  logic   [   5:0] regs$dump_out$017;
  logic   [   5:0] regs$dump_out$018;
  logic   [   5:0] regs$dump_out$019;
  logic   [   5:0] regs$dump_out$020;
  logic   [   5:0] regs$dump_out$021;
  logic   [   5:0] regs$dump_out$022;
  logic   [   5:0] regs$dump_out$023;
  logic   [   5:0] regs$dump_out$024;
  logic   [   5:0] regs$dump_out$025;
  logic   [   5:0] regs$dump_out$026;
  logic   [   5:0] regs$dump_out$027;
  logic   [   5:0] regs$dump_out$028;
  logic   [   5:0] regs$dump_out$029;
  logic   [   5:0] regs$dump_out$030;
  logic   [   5:0] regs$dump_out$031;

  RegisterFile_0x7c767f76bd64c12c regs
  (
    .set_in_$000    ( regs$set_in_$000 ),
    .set_in_$001    ( regs$set_in_$001 ),
    .set_in_$002    ( regs$set_in_$002 ),
    .set_in_$003    ( regs$set_in_$003 ),
    .set_in_$004    ( regs$set_in_$004 ),
    .set_in_$005    ( regs$set_in_$005 ),
    .set_in_$006    ( regs$set_in_$006 ),
    .set_in_$007    ( regs$set_in_$007 ),
    .set_in_$008    ( regs$set_in_$008 ),
    .set_in_$009    ( regs$set_in_$009 ),
    .set_in_$010    ( regs$set_in_$010 ),
    .set_in_$011    ( regs$set_in_$011 ),
    .set_in_$012    ( regs$set_in_$012 ),
    .set_in_$013    ( regs$set_in_$013 ),
    .set_in_$014    ( regs$set_in_$014 ),
    .set_in_$015    ( regs$set_in_$015 ),
    .set_in_$016    ( regs$set_in_$016 ),
    .set_in_$017    ( regs$set_in_$017 ),
    .set_in_$018    ( regs$set_in_$018 ),
    .set_in_$019    ( regs$set_in_$019 ),
    .set_in_$020    ( regs$set_in_$020 ),
    .set_in_$021    ( regs$set_in_$021 ),
    .set_in_$022    ( regs$set_in_$022 ),
    .set_in_$023    ( regs$set_in_$023 ),
    .set_in_$024    ( regs$set_in_$024 ),
    .set_in_$025    ( regs$set_in_$025 ),
    .set_in_$026    ( regs$set_in_$026 ),
    .set_in_$027    ( regs$set_in_$027 ),
    .set_in_$028    ( regs$set_in_$028 ),
    .set_in_$029    ( regs$set_in_$029 ),
    .set_in_$030    ( regs$set_in_$030 ),
    .set_in_$031    ( regs$set_in_$031 ),
    .set_call       ( regs$set_call ),
    .clk            ( regs$clk ),
    .write_addr$000 ( regs$write_addr$000 ),
    .read_addr$000  ( regs$read_addr$000 ),
    .read_addr$001  ( regs$read_addr$001 ),
    .write_call$000 ( regs$write_call$000 ),
    .write_data$000 ( regs$write_data$000 ),
    .reset          ( regs$reset ),
    .read_data$000  ( regs$read_data$000 ),
    .read_data$001  ( regs$read_data$001 ),
    .dump_out$000   ( regs$dump_out$000 ),
    .dump_out$001   ( regs$dump_out$001 ),
    .dump_out$002   ( regs$dump_out$002 ),
    .dump_out$003   ( regs$dump_out$003 ),
    .dump_out$004   ( regs$dump_out$004 ),
    .dump_out$005   ( regs$dump_out$005 ),
    .dump_out$006   ( regs$dump_out$006 ),
    .dump_out$007   ( regs$dump_out$007 ),
    .dump_out$008   ( regs$dump_out$008 ),
    .dump_out$009   ( regs$dump_out$009 ),
    .dump_out$010   ( regs$dump_out$010 ),
    .dump_out$011   ( regs$dump_out$011 ),
    .dump_out$012   ( regs$dump_out$012 ),
    .dump_out$013   ( regs$dump_out$013 ),
    .dump_out$014   ( regs$dump_out$014 ),
    .dump_out$015   ( regs$dump_out$015 ),
    .dump_out$016   ( regs$dump_out$016 ),
    .dump_out$017   ( regs$dump_out$017 ),
    .dump_out$018   ( regs$dump_out$018 ),
    .dump_out$019   ( regs$dump_out$019 ),
    .dump_out$020   ( regs$dump_out$020 ),
    .dump_out$021   ( regs$dump_out$021 ),
    .dump_out$022   ( regs$dump_out$022 ),
    .dump_out$023   ( regs$dump_out$023 ),
    .dump_out$024   ( regs$dump_out$024 ),
    .dump_out$025   ( regs$dump_out$025 ),
    .dump_out$026   ( regs$dump_out$026 ),
    .dump_out$027   ( regs$dump_out$027 ),
    .dump_out$028   ( regs$dump_out$028 ),
    .dump_out$029   ( regs$dump_out$029 ),
    .dump_out$030   ( regs$dump_out$030 ),
    .dump_out$031   ( regs$dump_out$031 )
  );

  // snapshot_muxes$000 temporaries
  logic   [   5:0] snapshot_muxes$000$mux_in_$000;
  logic   [   5:0] snapshot_muxes$000$mux_in_$001;
  logic   [   0:0] snapshot_muxes$000$clk;
  logic   [   0:0] snapshot_muxes$000$reset;
  logic   [   0:0] snapshot_muxes$000$mux_select;
  logic   [   5:0] snapshot_muxes$000$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$000
  (
    .mux_in_$000 ( snapshot_muxes$000$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$000$mux_in_$001 ),
    .clk         ( snapshot_muxes$000$clk ),
    .reset       ( snapshot_muxes$000$reset ),
    .mux_select  ( snapshot_muxes$000$mux_select ),
    .mux_out     ( snapshot_muxes$000$mux_out )
  );

  // snapshot_muxes$001 temporaries
  logic   [   5:0] snapshot_muxes$001$mux_in_$000;
  logic   [   5:0] snapshot_muxes$001$mux_in_$001;
  logic   [   0:0] snapshot_muxes$001$clk;
  logic   [   0:0] snapshot_muxes$001$reset;
  logic   [   0:0] snapshot_muxes$001$mux_select;
  logic   [   5:0] snapshot_muxes$001$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$001
  (
    .mux_in_$000 ( snapshot_muxes$001$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$001$mux_in_$001 ),
    .clk         ( snapshot_muxes$001$clk ),
    .reset       ( snapshot_muxes$001$reset ),
    .mux_select  ( snapshot_muxes$001$mux_select ),
    .mux_out     ( snapshot_muxes$001$mux_out )
  );

  // snapshot_muxes$002 temporaries
  logic   [   5:0] snapshot_muxes$002$mux_in_$000;
  logic   [   5:0] snapshot_muxes$002$mux_in_$001;
  logic   [   0:0] snapshot_muxes$002$clk;
  logic   [   0:0] snapshot_muxes$002$reset;
  logic   [   0:0] snapshot_muxes$002$mux_select;
  logic   [   5:0] snapshot_muxes$002$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$002
  (
    .mux_in_$000 ( snapshot_muxes$002$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$002$mux_in_$001 ),
    .clk         ( snapshot_muxes$002$clk ),
    .reset       ( snapshot_muxes$002$reset ),
    .mux_select  ( snapshot_muxes$002$mux_select ),
    .mux_out     ( snapshot_muxes$002$mux_out )
  );

  // snapshot_muxes$003 temporaries
  logic   [   5:0] snapshot_muxes$003$mux_in_$000;
  logic   [   5:0] snapshot_muxes$003$mux_in_$001;
  logic   [   0:0] snapshot_muxes$003$clk;
  logic   [   0:0] snapshot_muxes$003$reset;
  logic   [   0:0] snapshot_muxes$003$mux_select;
  logic   [   5:0] snapshot_muxes$003$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$003
  (
    .mux_in_$000 ( snapshot_muxes$003$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$003$mux_in_$001 ),
    .clk         ( snapshot_muxes$003$clk ),
    .reset       ( snapshot_muxes$003$reset ),
    .mux_select  ( snapshot_muxes$003$mux_select ),
    .mux_out     ( snapshot_muxes$003$mux_out )
  );

  // snapshot_muxes$004 temporaries
  logic   [   5:0] snapshot_muxes$004$mux_in_$000;
  logic   [   5:0] snapshot_muxes$004$mux_in_$001;
  logic   [   0:0] snapshot_muxes$004$clk;
  logic   [   0:0] snapshot_muxes$004$reset;
  logic   [   0:0] snapshot_muxes$004$mux_select;
  logic   [   5:0] snapshot_muxes$004$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$004
  (
    .mux_in_$000 ( snapshot_muxes$004$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$004$mux_in_$001 ),
    .clk         ( snapshot_muxes$004$clk ),
    .reset       ( snapshot_muxes$004$reset ),
    .mux_select  ( snapshot_muxes$004$mux_select ),
    .mux_out     ( snapshot_muxes$004$mux_out )
  );

  // snapshot_muxes$005 temporaries
  logic   [   5:0] snapshot_muxes$005$mux_in_$000;
  logic   [   5:0] snapshot_muxes$005$mux_in_$001;
  logic   [   0:0] snapshot_muxes$005$clk;
  logic   [   0:0] snapshot_muxes$005$reset;
  logic   [   0:0] snapshot_muxes$005$mux_select;
  logic   [   5:0] snapshot_muxes$005$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$005
  (
    .mux_in_$000 ( snapshot_muxes$005$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$005$mux_in_$001 ),
    .clk         ( snapshot_muxes$005$clk ),
    .reset       ( snapshot_muxes$005$reset ),
    .mux_select  ( snapshot_muxes$005$mux_select ),
    .mux_out     ( snapshot_muxes$005$mux_out )
  );

  // snapshot_muxes$006 temporaries
  logic   [   5:0] snapshot_muxes$006$mux_in_$000;
  logic   [   5:0] snapshot_muxes$006$mux_in_$001;
  logic   [   0:0] snapshot_muxes$006$clk;
  logic   [   0:0] snapshot_muxes$006$reset;
  logic   [   0:0] snapshot_muxes$006$mux_select;
  logic   [   5:0] snapshot_muxes$006$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$006
  (
    .mux_in_$000 ( snapshot_muxes$006$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$006$mux_in_$001 ),
    .clk         ( snapshot_muxes$006$clk ),
    .reset       ( snapshot_muxes$006$reset ),
    .mux_select  ( snapshot_muxes$006$mux_select ),
    .mux_out     ( snapshot_muxes$006$mux_out )
  );

  // snapshot_muxes$007 temporaries
  logic   [   5:0] snapshot_muxes$007$mux_in_$000;
  logic   [   5:0] snapshot_muxes$007$mux_in_$001;
  logic   [   0:0] snapshot_muxes$007$clk;
  logic   [   0:0] snapshot_muxes$007$reset;
  logic   [   0:0] snapshot_muxes$007$mux_select;
  logic   [   5:0] snapshot_muxes$007$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$007
  (
    .mux_in_$000 ( snapshot_muxes$007$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$007$mux_in_$001 ),
    .clk         ( snapshot_muxes$007$clk ),
    .reset       ( snapshot_muxes$007$reset ),
    .mux_select  ( snapshot_muxes$007$mux_select ),
    .mux_out     ( snapshot_muxes$007$mux_out )
  );

  // snapshot_muxes$008 temporaries
  logic   [   5:0] snapshot_muxes$008$mux_in_$000;
  logic   [   5:0] snapshot_muxes$008$mux_in_$001;
  logic   [   0:0] snapshot_muxes$008$clk;
  logic   [   0:0] snapshot_muxes$008$reset;
  logic   [   0:0] snapshot_muxes$008$mux_select;
  logic   [   5:0] snapshot_muxes$008$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$008
  (
    .mux_in_$000 ( snapshot_muxes$008$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$008$mux_in_$001 ),
    .clk         ( snapshot_muxes$008$clk ),
    .reset       ( snapshot_muxes$008$reset ),
    .mux_select  ( snapshot_muxes$008$mux_select ),
    .mux_out     ( snapshot_muxes$008$mux_out )
  );

  // snapshot_muxes$009 temporaries
  logic   [   5:0] snapshot_muxes$009$mux_in_$000;
  logic   [   5:0] snapshot_muxes$009$mux_in_$001;
  logic   [   0:0] snapshot_muxes$009$clk;
  logic   [   0:0] snapshot_muxes$009$reset;
  logic   [   0:0] snapshot_muxes$009$mux_select;
  logic   [   5:0] snapshot_muxes$009$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$009
  (
    .mux_in_$000 ( snapshot_muxes$009$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$009$mux_in_$001 ),
    .clk         ( snapshot_muxes$009$clk ),
    .reset       ( snapshot_muxes$009$reset ),
    .mux_select  ( snapshot_muxes$009$mux_select ),
    .mux_out     ( snapshot_muxes$009$mux_out )
  );

  // snapshot_muxes$010 temporaries
  logic   [   5:0] snapshot_muxes$010$mux_in_$000;
  logic   [   5:0] snapshot_muxes$010$mux_in_$001;
  logic   [   0:0] snapshot_muxes$010$clk;
  logic   [   0:0] snapshot_muxes$010$reset;
  logic   [   0:0] snapshot_muxes$010$mux_select;
  logic   [   5:0] snapshot_muxes$010$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$010
  (
    .mux_in_$000 ( snapshot_muxes$010$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$010$mux_in_$001 ),
    .clk         ( snapshot_muxes$010$clk ),
    .reset       ( snapshot_muxes$010$reset ),
    .mux_select  ( snapshot_muxes$010$mux_select ),
    .mux_out     ( snapshot_muxes$010$mux_out )
  );

  // snapshot_muxes$011 temporaries
  logic   [   5:0] snapshot_muxes$011$mux_in_$000;
  logic   [   5:0] snapshot_muxes$011$mux_in_$001;
  logic   [   0:0] snapshot_muxes$011$clk;
  logic   [   0:0] snapshot_muxes$011$reset;
  logic   [   0:0] snapshot_muxes$011$mux_select;
  logic   [   5:0] snapshot_muxes$011$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$011
  (
    .mux_in_$000 ( snapshot_muxes$011$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$011$mux_in_$001 ),
    .clk         ( snapshot_muxes$011$clk ),
    .reset       ( snapshot_muxes$011$reset ),
    .mux_select  ( snapshot_muxes$011$mux_select ),
    .mux_out     ( snapshot_muxes$011$mux_out )
  );

  // snapshot_muxes$012 temporaries
  logic   [   5:0] snapshot_muxes$012$mux_in_$000;
  logic   [   5:0] snapshot_muxes$012$mux_in_$001;
  logic   [   0:0] snapshot_muxes$012$clk;
  logic   [   0:0] snapshot_muxes$012$reset;
  logic   [   0:0] snapshot_muxes$012$mux_select;
  logic   [   5:0] snapshot_muxes$012$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$012
  (
    .mux_in_$000 ( snapshot_muxes$012$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$012$mux_in_$001 ),
    .clk         ( snapshot_muxes$012$clk ),
    .reset       ( snapshot_muxes$012$reset ),
    .mux_select  ( snapshot_muxes$012$mux_select ),
    .mux_out     ( snapshot_muxes$012$mux_out )
  );

  // snapshot_muxes$013 temporaries
  logic   [   5:0] snapshot_muxes$013$mux_in_$000;
  logic   [   5:0] snapshot_muxes$013$mux_in_$001;
  logic   [   0:0] snapshot_muxes$013$clk;
  logic   [   0:0] snapshot_muxes$013$reset;
  logic   [   0:0] snapshot_muxes$013$mux_select;
  logic   [   5:0] snapshot_muxes$013$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$013
  (
    .mux_in_$000 ( snapshot_muxes$013$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$013$mux_in_$001 ),
    .clk         ( snapshot_muxes$013$clk ),
    .reset       ( snapshot_muxes$013$reset ),
    .mux_select  ( snapshot_muxes$013$mux_select ),
    .mux_out     ( snapshot_muxes$013$mux_out )
  );

  // snapshot_muxes$014 temporaries
  logic   [   5:0] snapshot_muxes$014$mux_in_$000;
  logic   [   5:0] snapshot_muxes$014$mux_in_$001;
  logic   [   0:0] snapshot_muxes$014$clk;
  logic   [   0:0] snapshot_muxes$014$reset;
  logic   [   0:0] snapshot_muxes$014$mux_select;
  logic   [   5:0] snapshot_muxes$014$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$014
  (
    .mux_in_$000 ( snapshot_muxes$014$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$014$mux_in_$001 ),
    .clk         ( snapshot_muxes$014$clk ),
    .reset       ( snapshot_muxes$014$reset ),
    .mux_select  ( snapshot_muxes$014$mux_select ),
    .mux_out     ( snapshot_muxes$014$mux_out )
  );

  // snapshot_muxes$015 temporaries
  logic   [   5:0] snapshot_muxes$015$mux_in_$000;
  logic   [   5:0] snapshot_muxes$015$mux_in_$001;
  logic   [   0:0] snapshot_muxes$015$clk;
  logic   [   0:0] snapshot_muxes$015$reset;
  logic   [   0:0] snapshot_muxes$015$mux_select;
  logic   [   5:0] snapshot_muxes$015$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$015
  (
    .mux_in_$000 ( snapshot_muxes$015$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$015$mux_in_$001 ),
    .clk         ( snapshot_muxes$015$clk ),
    .reset       ( snapshot_muxes$015$reset ),
    .mux_select  ( snapshot_muxes$015$mux_select ),
    .mux_out     ( snapshot_muxes$015$mux_out )
  );

  // snapshot_muxes$016 temporaries
  logic   [   5:0] snapshot_muxes$016$mux_in_$000;
  logic   [   5:0] snapshot_muxes$016$mux_in_$001;
  logic   [   0:0] snapshot_muxes$016$clk;
  logic   [   0:0] snapshot_muxes$016$reset;
  logic   [   0:0] snapshot_muxes$016$mux_select;
  logic   [   5:0] snapshot_muxes$016$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$016
  (
    .mux_in_$000 ( snapshot_muxes$016$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$016$mux_in_$001 ),
    .clk         ( snapshot_muxes$016$clk ),
    .reset       ( snapshot_muxes$016$reset ),
    .mux_select  ( snapshot_muxes$016$mux_select ),
    .mux_out     ( snapshot_muxes$016$mux_out )
  );

  // snapshot_muxes$017 temporaries
  logic   [   5:0] snapshot_muxes$017$mux_in_$000;
  logic   [   5:0] snapshot_muxes$017$mux_in_$001;
  logic   [   0:0] snapshot_muxes$017$clk;
  logic   [   0:0] snapshot_muxes$017$reset;
  logic   [   0:0] snapshot_muxes$017$mux_select;
  logic   [   5:0] snapshot_muxes$017$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$017
  (
    .mux_in_$000 ( snapshot_muxes$017$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$017$mux_in_$001 ),
    .clk         ( snapshot_muxes$017$clk ),
    .reset       ( snapshot_muxes$017$reset ),
    .mux_select  ( snapshot_muxes$017$mux_select ),
    .mux_out     ( snapshot_muxes$017$mux_out )
  );

  // snapshot_muxes$018 temporaries
  logic   [   5:0] snapshot_muxes$018$mux_in_$000;
  logic   [   5:0] snapshot_muxes$018$mux_in_$001;
  logic   [   0:0] snapshot_muxes$018$clk;
  logic   [   0:0] snapshot_muxes$018$reset;
  logic   [   0:0] snapshot_muxes$018$mux_select;
  logic   [   5:0] snapshot_muxes$018$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$018
  (
    .mux_in_$000 ( snapshot_muxes$018$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$018$mux_in_$001 ),
    .clk         ( snapshot_muxes$018$clk ),
    .reset       ( snapshot_muxes$018$reset ),
    .mux_select  ( snapshot_muxes$018$mux_select ),
    .mux_out     ( snapshot_muxes$018$mux_out )
  );

  // snapshot_muxes$019 temporaries
  logic   [   5:0] snapshot_muxes$019$mux_in_$000;
  logic   [   5:0] snapshot_muxes$019$mux_in_$001;
  logic   [   0:0] snapshot_muxes$019$clk;
  logic   [   0:0] snapshot_muxes$019$reset;
  logic   [   0:0] snapshot_muxes$019$mux_select;
  logic   [   5:0] snapshot_muxes$019$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$019
  (
    .mux_in_$000 ( snapshot_muxes$019$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$019$mux_in_$001 ),
    .clk         ( snapshot_muxes$019$clk ),
    .reset       ( snapshot_muxes$019$reset ),
    .mux_select  ( snapshot_muxes$019$mux_select ),
    .mux_out     ( snapshot_muxes$019$mux_out )
  );

  // snapshot_muxes$020 temporaries
  logic   [   5:0] snapshot_muxes$020$mux_in_$000;
  logic   [   5:0] snapshot_muxes$020$mux_in_$001;
  logic   [   0:0] snapshot_muxes$020$clk;
  logic   [   0:0] snapshot_muxes$020$reset;
  logic   [   0:0] snapshot_muxes$020$mux_select;
  logic   [   5:0] snapshot_muxes$020$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$020
  (
    .mux_in_$000 ( snapshot_muxes$020$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$020$mux_in_$001 ),
    .clk         ( snapshot_muxes$020$clk ),
    .reset       ( snapshot_muxes$020$reset ),
    .mux_select  ( snapshot_muxes$020$mux_select ),
    .mux_out     ( snapshot_muxes$020$mux_out )
  );

  // snapshot_muxes$021 temporaries
  logic   [   5:0] snapshot_muxes$021$mux_in_$000;
  logic   [   5:0] snapshot_muxes$021$mux_in_$001;
  logic   [   0:0] snapshot_muxes$021$clk;
  logic   [   0:0] snapshot_muxes$021$reset;
  logic   [   0:0] snapshot_muxes$021$mux_select;
  logic   [   5:0] snapshot_muxes$021$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$021
  (
    .mux_in_$000 ( snapshot_muxes$021$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$021$mux_in_$001 ),
    .clk         ( snapshot_muxes$021$clk ),
    .reset       ( snapshot_muxes$021$reset ),
    .mux_select  ( snapshot_muxes$021$mux_select ),
    .mux_out     ( snapshot_muxes$021$mux_out )
  );

  // snapshot_muxes$022 temporaries
  logic   [   5:0] snapshot_muxes$022$mux_in_$000;
  logic   [   5:0] snapshot_muxes$022$mux_in_$001;
  logic   [   0:0] snapshot_muxes$022$clk;
  logic   [   0:0] snapshot_muxes$022$reset;
  logic   [   0:0] snapshot_muxes$022$mux_select;
  logic   [   5:0] snapshot_muxes$022$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$022
  (
    .mux_in_$000 ( snapshot_muxes$022$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$022$mux_in_$001 ),
    .clk         ( snapshot_muxes$022$clk ),
    .reset       ( snapshot_muxes$022$reset ),
    .mux_select  ( snapshot_muxes$022$mux_select ),
    .mux_out     ( snapshot_muxes$022$mux_out )
  );

  // snapshot_muxes$023 temporaries
  logic   [   5:0] snapshot_muxes$023$mux_in_$000;
  logic   [   5:0] snapshot_muxes$023$mux_in_$001;
  logic   [   0:0] snapshot_muxes$023$clk;
  logic   [   0:0] snapshot_muxes$023$reset;
  logic   [   0:0] snapshot_muxes$023$mux_select;
  logic   [   5:0] snapshot_muxes$023$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$023
  (
    .mux_in_$000 ( snapshot_muxes$023$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$023$mux_in_$001 ),
    .clk         ( snapshot_muxes$023$clk ),
    .reset       ( snapshot_muxes$023$reset ),
    .mux_select  ( snapshot_muxes$023$mux_select ),
    .mux_out     ( snapshot_muxes$023$mux_out )
  );

  // snapshot_muxes$024 temporaries
  logic   [   5:0] snapshot_muxes$024$mux_in_$000;
  logic   [   5:0] snapshot_muxes$024$mux_in_$001;
  logic   [   0:0] snapshot_muxes$024$clk;
  logic   [   0:0] snapshot_muxes$024$reset;
  logic   [   0:0] snapshot_muxes$024$mux_select;
  logic   [   5:0] snapshot_muxes$024$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$024
  (
    .mux_in_$000 ( snapshot_muxes$024$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$024$mux_in_$001 ),
    .clk         ( snapshot_muxes$024$clk ),
    .reset       ( snapshot_muxes$024$reset ),
    .mux_select  ( snapshot_muxes$024$mux_select ),
    .mux_out     ( snapshot_muxes$024$mux_out )
  );

  // snapshot_muxes$025 temporaries
  logic   [   5:0] snapshot_muxes$025$mux_in_$000;
  logic   [   5:0] snapshot_muxes$025$mux_in_$001;
  logic   [   0:0] snapshot_muxes$025$clk;
  logic   [   0:0] snapshot_muxes$025$reset;
  logic   [   0:0] snapshot_muxes$025$mux_select;
  logic   [   5:0] snapshot_muxes$025$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$025
  (
    .mux_in_$000 ( snapshot_muxes$025$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$025$mux_in_$001 ),
    .clk         ( snapshot_muxes$025$clk ),
    .reset       ( snapshot_muxes$025$reset ),
    .mux_select  ( snapshot_muxes$025$mux_select ),
    .mux_out     ( snapshot_muxes$025$mux_out )
  );

  // snapshot_muxes$026 temporaries
  logic   [   5:0] snapshot_muxes$026$mux_in_$000;
  logic   [   5:0] snapshot_muxes$026$mux_in_$001;
  logic   [   0:0] snapshot_muxes$026$clk;
  logic   [   0:0] snapshot_muxes$026$reset;
  logic   [   0:0] snapshot_muxes$026$mux_select;
  logic   [   5:0] snapshot_muxes$026$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$026
  (
    .mux_in_$000 ( snapshot_muxes$026$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$026$mux_in_$001 ),
    .clk         ( snapshot_muxes$026$clk ),
    .reset       ( snapshot_muxes$026$reset ),
    .mux_select  ( snapshot_muxes$026$mux_select ),
    .mux_out     ( snapshot_muxes$026$mux_out )
  );

  // snapshot_muxes$027 temporaries
  logic   [   5:0] snapshot_muxes$027$mux_in_$000;
  logic   [   5:0] snapshot_muxes$027$mux_in_$001;
  logic   [   0:0] snapshot_muxes$027$clk;
  logic   [   0:0] snapshot_muxes$027$reset;
  logic   [   0:0] snapshot_muxes$027$mux_select;
  logic   [   5:0] snapshot_muxes$027$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$027
  (
    .mux_in_$000 ( snapshot_muxes$027$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$027$mux_in_$001 ),
    .clk         ( snapshot_muxes$027$clk ),
    .reset       ( snapshot_muxes$027$reset ),
    .mux_select  ( snapshot_muxes$027$mux_select ),
    .mux_out     ( snapshot_muxes$027$mux_out )
  );

  // snapshot_muxes$028 temporaries
  logic   [   5:0] snapshot_muxes$028$mux_in_$000;
  logic   [   5:0] snapshot_muxes$028$mux_in_$001;
  logic   [   0:0] snapshot_muxes$028$clk;
  logic   [   0:0] snapshot_muxes$028$reset;
  logic   [   0:0] snapshot_muxes$028$mux_select;
  logic   [   5:0] snapshot_muxes$028$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$028
  (
    .mux_in_$000 ( snapshot_muxes$028$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$028$mux_in_$001 ),
    .clk         ( snapshot_muxes$028$clk ),
    .reset       ( snapshot_muxes$028$reset ),
    .mux_select  ( snapshot_muxes$028$mux_select ),
    .mux_out     ( snapshot_muxes$028$mux_out )
  );

  // snapshot_muxes$029 temporaries
  logic   [   5:0] snapshot_muxes$029$mux_in_$000;
  logic   [   5:0] snapshot_muxes$029$mux_in_$001;
  logic   [   0:0] snapshot_muxes$029$clk;
  logic   [   0:0] snapshot_muxes$029$reset;
  logic   [   0:0] snapshot_muxes$029$mux_select;
  logic   [   5:0] snapshot_muxes$029$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$029
  (
    .mux_in_$000 ( snapshot_muxes$029$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$029$mux_in_$001 ),
    .clk         ( snapshot_muxes$029$clk ),
    .reset       ( snapshot_muxes$029$reset ),
    .mux_select  ( snapshot_muxes$029$mux_select ),
    .mux_out     ( snapshot_muxes$029$mux_out )
  );

  // snapshot_muxes$030 temporaries
  logic   [   5:0] snapshot_muxes$030$mux_in_$000;
  logic   [   5:0] snapshot_muxes$030$mux_in_$001;
  logic   [   0:0] snapshot_muxes$030$clk;
  logic   [   0:0] snapshot_muxes$030$reset;
  logic   [   0:0] snapshot_muxes$030$mux_select;
  logic   [   5:0] snapshot_muxes$030$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$030
  (
    .mux_in_$000 ( snapshot_muxes$030$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$030$mux_in_$001 ),
    .clk         ( snapshot_muxes$030$clk ),
    .reset       ( snapshot_muxes$030$reset ),
    .mux_select  ( snapshot_muxes$030$mux_select ),
    .mux_out     ( snapshot_muxes$030$mux_out )
  );

  // snapshot_muxes$031 temporaries
  logic   [   5:0] snapshot_muxes$031$mux_in_$000;
  logic   [   5:0] snapshot_muxes$031$mux_in_$001;
  logic   [   0:0] snapshot_muxes$031$clk;
  logic   [   0:0] snapshot_muxes$031$reset;
  logic   [   0:0] snapshot_muxes$031$mux_select;
  logic   [   5:0] snapshot_muxes$031$mux_out;

  Mux_0x387678144da2c8e snapshot_muxes$031
  (
    .mux_in_$000 ( snapshot_muxes$031$mux_in_$000 ),
    .mux_in_$001 ( snapshot_muxes$031$mux_in_$001 ),
    .clk         ( snapshot_muxes$031$clk ),
    .reset       ( snapshot_muxes$031$reset ),
    .mux_select  ( snapshot_muxes$031$mux_select ),
    .mux_out     ( snapshot_muxes$031$mux_out )
  );

  // set_muxes$000 temporaries
  logic   [   5:0] set_muxes$000$mux_in_$000;
  logic   [   5:0] set_muxes$000$mux_in_$001;
  logic   [   0:0] set_muxes$000$clk;
  logic   [   0:0] set_muxes$000$reset;
  logic   [   0:0] set_muxes$000$mux_select;
  logic   [   5:0] set_muxes$000$mux_out;

  Mux_0x387678144da2c8e set_muxes$000
  (
    .mux_in_$000 ( set_muxes$000$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$000$mux_in_$001 ),
    .clk         ( set_muxes$000$clk ),
    .reset       ( set_muxes$000$reset ),
    .mux_select  ( set_muxes$000$mux_select ),
    .mux_out     ( set_muxes$000$mux_out )
  );

  // set_muxes$001 temporaries
  logic   [   5:0] set_muxes$001$mux_in_$000;
  logic   [   5:0] set_muxes$001$mux_in_$001;
  logic   [   0:0] set_muxes$001$clk;
  logic   [   0:0] set_muxes$001$reset;
  logic   [   0:0] set_muxes$001$mux_select;
  logic   [   5:0] set_muxes$001$mux_out;

  Mux_0x387678144da2c8e set_muxes$001
  (
    .mux_in_$000 ( set_muxes$001$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$001$mux_in_$001 ),
    .clk         ( set_muxes$001$clk ),
    .reset       ( set_muxes$001$reset ),
    .mux_select  ( set_muxes$001$mux_select ),
    .mux_out     ( set_muxes$001$mux_out )
  );

  // set_muxes$002 temporaries
  logic   [   5:0] set_muxes$002$mux_in_$000;
  logic   [   5:0] set_muxes$002$mux_in_$001;
  logic   [   0:0] set_muxes$002$clk;
  logic   [   0:0] set_muxes$002$reset;
  logic   [   0:0] set_muxes$002$mux_select;
  logic   [   5:0] set_muxes$002$mux_out;

  Mux_0x387678144da2c8e set_muxes$002
  (
    .mux_in_$000 ( set_muxes$002$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$002$mux_in_$001 ),
    .clk         ( set_muxes$002$clk ),
    .reset       ( set_muxes$002$reset ),
    .mux_select  ( set_muxes$002$mux_select ),
    .mux_out     ( set_muxes$002$mux_out )
  );

  // set_muxes$003 temporaries
  logic   [   5:0] set_muxes$003$mux_in_$000;
  logic   [   5:0] set_muxes$003$mux_in_$001;
  logic   [   0:0] set_muxes$003$clk;
  logic   [   0:0] set_muxes$003$reset;
  logic   [   0:0] set_muxes$003$mux_select;
  logic   [   5:0] set_muxes$003$mux_out;

  Mux_0x387678144da2c8e set_muxes$003
  (
    .mux_in_$000 ( set_muxes$003$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$003$mux_in_$001 ),
    .clk         ( set_muxes$003$clk ),
    .reset       ( set_muxes$003$reset ),
    .mux_select  ( set_muxes$003$mux_select ),
    .mux_out     ( set_muxes$003$mux_out )
  );

  // set_muxes$004 temporaries
  logic   [   5:0] set_muxes$004$mux_in_$000;
  logic   [   5:0] set_muxes$004$mux_in_$001;
  logic   [   0:0] set_muxes$004$clk;
  logic   [   0:0] set_muxes$004$reset;
  logic   [   0:0] set_muxes$004$mux_select;
  logic   [   5:0] set_muxes$004$mux_out;

  Mux_0x387678144da2c8e set_muxes$004
  (
    .mux_in_$000 ( set_muxes$004$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$004$mux_in_$001 ),
    .clk         ( set_muxes$004$clk ),
    .reset       ( set_muxes$004$reset ),
    .mux_select  ( set_muxes$004$mux_select ),
    .mux_out     ( set_muxes$004$mux_out )
  );

  // set_muxes$005 temporaries
  logic   [   5:0] set_muxes$005$mux_in_$000;
  logic   [   5:0] set_muxes$005$mux_in_$001;
  logic   [   0:0] set_muxes$005$clk;
  logic   [   0:0] set_muxes$005$reset;
  logic   [   0:0] set_muxes$005$mux_select;
  logic   [   5:0] set_muxes$005$mux_out;

  Mux_0x387678144da2c8e set_muxes$005
  (
    .mux_in_$000 ( set_muxes$005$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$005$mux_in_$001 ),
    .clk         ( set_muxes$005$clk ),
    .reset       ( set_muxes$005$reset ),
    .mux_select  ( set_muxes$005$mux_select ),
    .mux_out     ( set_muxes$005$mux_out )
  );

  // set_muxes$006 temporaries
  logic   [   5:0] set_muxes$006$mux_in_$000;
  logic   [   5:0] set_muxes$006$mux_in_$001;
  logic   [   0:0] set_muxes$006$clk;
  logic   [   0:0] set_muxes$006$reset;
  logic   [   0:0] set_muxes$006$mux_select;
  logic   [   5:0] set_muxes$006$mux_out;

  Mux_0x387678144da2c8e set_muxes$006
  (
    .mux_in_$000 ( set_muxes$006$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$006$mux_in_$001 ),
    .clk         ( set_muxes$006$clk ),
    .reset       ( set_muxes$006$reset ),
    .mux_select  ( set_muxes$006$mux_select ),
    .mux_out     ( set_muxes$006$mux_out )
  );

  // set_muxes$007 temporaries
  logic   [   5:0] set_muxes$007$mux_in_$000;
  logic   [   5:0] set_muxes$007$mux_in_$001;
  logic   [   0:0] set_muxes$007$clk;
  logic   [   0:0] set_muxes$007$reset;
  logic   [   0:0] set_muxes$007$mux_select;
  logic   [   5:0] set_muxes$007$mux_out;

  Mux_0x387678144da2c8e set_muxes$007
  (
    .mux_in_$000 ( set_muxes$007$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$007$mux_in_$001 ),
    .clk         ( set_muxes$007$clk ),
    .reset       ( set_muxes$007$reset ),
    .mux_select  ( set_muxes$007$mux_select ),
    .mux_out     ( set_muxes$007$mux_out )
  );

  // set_muxes$008 temporaries
  logic   [   5:0] set_muxes$008$mux_in_$000;
  logic   [   5:0] set_muxes$008$mux_in_$001;
  logic   [   0:0] set_muxes$008$clk;
  logic   [   0:0] set_muxes$008$reset;
  logic   [   0:0] set_muxes$008$mux_select;
  logic   [   5:0] set_muxes$008$mux_out;

  Mux_0x387678144da2c8e set_muxes$008
  (
    .mux_in_$000 ( set_muxes$008$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$008$mux_in_$001 ),
    .clk         ( set_muxes$008$clk ),
    .reset       ( set_muxes$008$reset ),
    .mux_select  ( set_muxes$008$mux_select ),
    .mux_out     ( set_muxes$008$mux_out )
  );

  // set_muxes$009 temporaries
  logic   [   5:0] set_muxes$009$mux_in_$000;
  logic   [   5:0] set_muxes$009$mux_in_$001;
  logic   [   0:0] set_muxes$009$clk;
  logic   [   0:0] set_muxes$009$reset;
  logic   [   0:0] set_muxes$009$mux_select;
  logic   [   5:0] set_muxes$009$mux_out;

  Mux_0x387678144da2c8e set_muxes$009
  (
    .mux_in_$000 ( set_muxes$009$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$009$mux_in_$001 ),
    .clk         ( set_muxes$009$clk ),
    .reset       ( set_muxes$009$reset ),
    .mux_select  ( set_muxes$009$mux_select ),
    .mux_out     ( set_muxes$009$mux_out )
  );

  // set_muxes$010 temporaries
  logic   [   5:0] set_muxes$010$mux_in_$000;
  logic   [   5:0] set_muxes$010$mux_in_$001;
  logic   [   0:0] set_muxes$010$clk;
  logic   [   0:0] set_muxes$010$reset;
  logic   [   0:0] set_muxes$010$mux_select;
  logic   [   5:0] set_muxes$010$mux_out;

  Mux_0x387678144da2c8e set_muxes$010
  (
    .mux_in_$000 ( set_muxes$010$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$010$mux_in_$001 ),
    .clk         ( set_muxes$010$clk ),
    .reset       ( set_muxes$010$reset ),
    .mux_select  ( set_muxes$010$mux_select ),
    .mux_out     ( set_muxes$010$mux_out )
  );

  // set_muxes$011 temporaries
  logic   [   5:0] set_muxes$011$mux_in_$000;
  logic   [   5:0] set_muxes$011$mux_in_$001;
  logic   [   0:0] set_muxes$011$clk;
  logic   [   0:0] set_muxes$011$reset;
  logic   [   0:0] set_muxes$011$mux_select;
  logic   [   5:0] set_muxes$011$mux_out;

  Mux_0x387678144da2c8e set_muxes$011
  (
    .mux_in_$000 ( set_muxes$011$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$011$mux_in_$001 ),
    .clk         ( set_muxes$011$clk ),
    .reset       ( set_muxes$011$reset ),
    .mux_select  ( set_muxes$011$mux_select ),
    .mux_out     ( set_muxes$011$mux_out )
  );

  // set_muxes$012 temporaries
  logic   [   5:0] set_muxes$012$mux_in_$000;
  logic   [   5:0] set_muxes$012$mux_in_$001;
  logic   [   0:0] set_muxes$012$clk;
  logic   [   0:0] set_muxes$012$reset;
  logic   [   0:0] set_muxes$012$mux_select;
  logic   [   5:0] set_muxes$012$mux_out;

  Mux_0x387678144da2c8e set_muxes$012
  (
    .mux_in_$000 ( set_muxes$012$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$012$mux_in_$001 ),
    .clk         ( set_muxes$012$clk ),
    .reset       ( set_muxes$012$reset ),
    .mux_select  ( set_muxes$012$mux_select ),
    .mux_out     ( set_muxes$012$mux_out )
  );

  // set_muxes$013 temporaries
  logic   [   5:0] set_muxes$013$mux_in_$000;
  logic   [   5:0] set_muxes$013$mux_in_$001;
  logic   [   0:0] set_muxes$013$clk;
  logic   [   0:0] set_muxes$013$reset;
  logic   [   0:0] set_muxes$013$mux_select;
  logic   [   5:0] set_muxes$013$mux_out;

  Mux_0x387678144da2c8e set_muxes$013
  (
    .mux_in_$000 ( set_muxes$013$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$013$mux_in_$001 ),
    .clk         ( set_muxes$013$clk ),
    .reset       ( set_muxes$013$reset ),
    .mux_select  ( set_muxes$013$mux_select ),
    .mux_out     ( set_muxes$013$mux_out )
  );

  // set_muxes$014 temporaries
  logic   [   5:0] set_muxes$014$mux_in_$000;
  logic   [   5:0] set_muxes$014$mux_in_$001;
  logic   [   0:0] set_muxes$014$clk;
  logic   [   0:0] set_muxes$014$reset;
  logic   [   0:0] set_muxes$014$mux_select;
  logic   [   5:0] set_muxes$014$mux_out;

  Mux_0x387678144da2c8e set_muxes$014
  (
    .mux_in_$000 ( set_muxes$014$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$014$mux_in_$001 ),
    .clk         ( set_muxes$014$clk ),
    .reset       ( set_muxes$014$reset ),
    .mux_select  ( set_muxes$014$mux_select ),
    .mux_out     ( set_muxes$014$mux_out )
  );

  // set_muxes$015 temporaries
  logic   [   5:0] set_muxes$015$mux_in_$000;
  logic   [   5:0] set_muxes$015$mux_in_$001;
  logic   [   0:0] set_muxes$015$clk;
  logic   [   0:0] set_muxes$015$reset;
  logic   [   0:0] set_muxes$015$mux_select;
  logic   [   5:0] set_muxes$015$mux_out;

  Mux_0x387678144da2c8e set_muxes$015
  (
    .mux_in_$000 ( set_muxes$015$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$015$mux_in_$001 ),
    .clk         ( set_muxes$015$clk ),
    .reset       ( set_muxes$015$reset ),
    .mux_select  ( set_muxes$015$mux_select ),
    .mux_out     ( set_muxes$015$mux_out )
  );

  // set_muxes$016 temporaries
  logic   [   5:0] set_muxes$016$mux_in_$000;
  logic   [   5:0] set_muxes$016$mux_in_$001;
  logic   [   0:0] set_muxes$016$clk;
  logic   [   0:0] set_muxes$016$reset;
  logic   [   0:0] set_muxes$016$mux_select;
  logic   [   5:0] set_muxes$016$mux_out;

  Mux_0x387678144da2c8e set_muxes$016
  (
    .mux_in_$000 ( set_muxes$016$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$016$mux_in_$001 ),
    .clk         ( set_muxes$016$clk ),
    .reset       ( set_muxes$016$reset ),
    .mux_select  ( set_muxes$016$mux_select ),
    .mux_out     ( set_muxes$016$mux_out )
  );

  // set_muxes$017 temporaries
  logic   [   5:0] set_muxes$017$mux_in_$000;
  logic   [   5:0] set_muxes$017$mux_in_$001;
  logic   [   0:0] set_muxes$017$clk;
  logic   [   0:0] set_muxes$017$reset;
  logic   [   0:0] set_muxes$017$mux_select;
  logic   [   5:0] set_muxes$017$mux_out;

  Mux_0x387678144da2c8e set_muxes$017
  (
    .mux_in_$000 ( set_muxes$017$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$017$mux_in_$001 ),
    .clk         ( set_muxes$017$clk ),
    .reset       ( set_muxes$017$reset ),
    .mux_select  ( set_muxes$017$mux_select ),
    .mux_out     ( set_muxes$017$mux_out )
  );

  // set_muxes$018 temporaries
  logic   [   5:0] set_muxes$018$mux_in_$000;
  logic   [   5:0] set_muxes$018$mux_in_$001;
  logic   [   0:0] set_muxes$018$clk;
  logic   [   0:0] set_muxes$018$reset;
  logic   [   0:0] set_muxes$018$mux_select;
  logic   [   5:0] set_muxes$018$mux_out;

  Mux_0x387678144da2c8e set_muxes$018
  (
    .mux_in_$000 ( set_muxes$018$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$018$mux_in_$001 ),
    .clk         ( set_muxes$018$clk ),
    .reset       ( set_muxes$018$reset ),
    .mux_select  ( set_muxes$018$mux_select ),
    .mux_out     ( set_muxes$018$mux_out )
  );

  // set_muxes$019 temporaries
  logic   [   5:0] set_muxes$019$mux_in_$000;
  logic   [   5:0] set_muxes$019$mux_in_$001;
  logic   [   0:0] set_muxes$019$clk;
  logic   [   0:0] set_muxes$019$reset;
  logic   [   0:0] set_muxes$019$mux_select;
  logic   [   5:0] set_muxes$019$mux_out;

  Mux_0x387678144da2c8e set_muxes$019
  (
    .mux_in_$000 ( set_muxes$019$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$019$mux_in_$001 ),
    .clk         ( set_muxes$019$clk ),
    .reset       ( set_muxes$019$reset ),
    .mux_select  ( set_muxes$019$mux_select ),
    .mux_out     ( set_muxes$019$mux_out )
  );

  // set_muxes$020 temporaries
  logic   [   5:0] set_muxes$020$mux_in_$000;
  logic   [   5:0] set_muxes$020$mux_in_$001;
  logic   [   0:0] set_muxes$020$clk;
  logic   [   0:0] set_muxes$020$reset;
  logic   [   0:0] set_muxes$020$mux_select;
  logic   [   5:0] set_muxes$020$mux_out;

  Mux_0x387678144da2c8e set_muxes$020
  (
    .mux_in_$000 ( set_muxes$020$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$020$mux_in_$001 ),
    .clk         ( set_muxes$020$clk ),
    .reset       ( set_muxes$020$reset ),
    .mux_select  ( set_muxes$020$mux_select ),
    .mux_out     ( set_muxes$020$mux_out )
  );

  // set_muxes$021 temporaries
  logic   [   5:0] set_muxes$021$mux_in_$000;
  logic   [   5:0] set_muxes$021$mux_in_$001;
  logic   [   0:0] set_muxes$021$clk;
  logic   [   0:0] set_muxes$021$reset;
  logic   [   0:0] set_muxes$021$mux_select;
  logic   [   5:0] set_muxes$021$mux_out;

  Mux_0x387678144da2c8e set_muxes$021
  (
    .mux_in_$000 ( set_muxes$021$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$021$mux_in_$001 ),
    .clk         ( set_muxes$021$clk ),
    .reset       ( set_muxes$021$reset ),
    .mux_select  ( set_muxes$021$mux_select ),
    .mux_out     ( set_muxes$021$mux_out )
  );

  // set_muxes$022 temporaries
  logic   [   5:0] set_muxes$022$mux_in_$000;
  logic   [   5:0] set_muxes$022$mux_in_$001;
  logic   [   0:0] set_muxes$022$clk;
  logic   [   0:0] set_muxes$022$reset;
  logic   [   0:0] set_muxes$022$mux_select;
  logic   [   5:0] set_muxes$022$mux_out;

  Mux_0x387678144da2c8e set_muxes$022
  (
    .mux_in_$000 ( set_muxes$022$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$022$mux_in_$001 ),
    .clk         ( set_muxes$022$clk ),
    .reset       ( set_muxes$022$reset ),
    .mux_select  ( set_muxes$022$mux_select ),
    .mux_out     ( set_muxes$022$mux_out )
  );

  // set_muxes$023 temporaries
  logic   [   5:0] set_muxes$023$mux_in_$000;
  logic   [   5:0] set_muxes$023$mux_in_$001;
  logic   [   0:0] set_muxes$023$clk;
  logic   [   0:0] set_muxes$023$reset;
  logic   [   0:0] set_muxes$023$mux_select;
  logic   [   5:0] set_muxes$023$mux_out;

  Mux_0x387678144da2c8e set_muxes$023
  (
    .mux_in_$000 ( set_muxes$023$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$023$mux_in_$001 ),
    .clk         ( set_muxes$023$clk ),
    .reset       ( set_muxes$023$reset ),
    .mux_select  ( set_muxes$023$mux_select ),
    .mux_out     ( set_muxes$023$mux_out )
  );

  // set_muxes$024 temporaries
  logic   [   5:0] set_muxes$024$mux_in_$000;
  logic   [   5:0] set_muxes$024$mux_in_$001;
  logic   [   0:0] set_muxes$024$clk;
  logic   [   0:0] set_muxes$024$reset;
  logic   [   0:0] set_muxes$024$mux_select;
  logic   [   5:0] set_muxes$024$mux_out;

  Mux_0x387678144da2c8e set_muxes$024
  (
    .mux_in_$000 ( set_muxes$024$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$024$mux_in_$001 ),
    .clk         ( set_muxes$024$clk ),
    .reset       ( set_muxes$024$reset ),
    .mux_select  ( set_muxes$024$mux_select ),
    .mux_out     ( set_muxes$024$mux_out )
  );

  // set_muxes$025 temporaries
  logic   [   5:0] set_muxes$025$mux_in_$000;
  logic   [   5:0] set_muxes$025$mux_in_$001;
  logic   [   0:0] set_muxes$025$clk;
  logic   [   0:0] set_muxes$025$reset;
  logic   [   0:0] set_muxes$025$mux_select;
  logic   [   5:0] set_muxes$025$mux_out;

  Mux_0x387678144da2c8e set_muxes$025
  (
    .mux_in_$000 ( set_muxes$025$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$025$mux_in_$001 ),
    .clk         ( set_muxes$025$clk ),
    .reset       ( set_muxes$025$reset ),
    .mux_select  ( set_muxes$025$mux_select ),
    .mux_out     ( set_muxes$025$mux_out )
  );

  // set_muxes$026 temporaries
  logic   [   5:0] set_muxes$026$mux_in_$000;
  logic   [   5:0] set_muxes$026$mux_in_$001;
  logic   [   0:0] set_muxes$026$clk;
  logic   [   0:0] set_muxes$026$reset;
  logic   [   0:0] set_muxes$026$mux_select;
  logic   [   5:0] set_muxes$026$mux_out;

  Mux_0x387678144da2c8e set_muxes$026
  (
    .mux_in_$000 ( set_muxes$026$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$026$mux_in_$001 ),
    .clk         ( set_muxes$026$clk ),
    .reset       ( set_muxes$026$reset ),
    .mux_select  ( set_muxes$026$mux_select ),
    .mux_out     ( set_muxes$026$mux_out )
  );

  // set_muxes$027 temporaries
  logic   [   5:0] set_muxes$027$mux_in_$000;
  logic   [   5:0] set_muxes$027$mux_in_$001;
  logic   [   0:0] set_muxes$027$clk;
  logic   [   0:0] set_muxes$027$reset;
  logic   [   0:0] set_muxes$027$mux_select;
  logic   [   5:0] set_muxes$027$mux_out;

  Mux_0x387678144da2c8e set_muxes$027
  (
    .mux_in_$000 ( set_muxes$027$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$027$mux_in_$001 ),
    .clk         ( set_muxes$027$clk ),
    .reset       ( set_muxes$027$reset ),
    .mux_select  ( set_muxes$027$mux_select ),
    .mux_out     ( set_muxes$027$mux_out )
  );

  // set_muxes$028 temporaries
  logic   [   5:0] set_muxes$028$mux_in_$000;
  logic   [   5:0] set_muxes$028$mux_in_$001;
  logic   [   0:0] set_muxes$028$clk;
  logic   [   0:0] set_muxes$028$reset;
  logic   [   0:0] set_muxes$028$mux_select;
  logic   [   5:0] set_muxes$028$mux_out;

  Mux_0x387678144da2c8e set_muxes$028
  (
    .mux_in_$000 ( set_muxes$028$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$028$mux_in_$001 ),
    .clk         ( set_muxes$028$clk ),
    .reset       ( set_muxes$028$reset ),
    .mux_select  ( set_muxes$028$mux_select ),
    .mux_out     ( set_muxes$028$mux_out )
  );

  // set_muxes$029 temporaries
  logic   [   5:0] set_muxes$029$mux_in_$000;
  logic   [   5:0] set_muxes$029$mux_in_$001;
  logic   [   0:0] set_muxes$029$clk;
  logic   [   0:0] set_muxes$029$reset;
  logic   [   0:0] set_muxes$029$mux_select;
  logic   [   5:0] set_muxes$029$mux_out;

  Mux_0x387678144da2c8e set_muxes$029
  (
    .mux_in_$000 ( set_muxes$029$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$029$mux_in_$001 ),
    .clk         ( set_muxes$029$clk ),
    .reset       ( set_muxes$029$reset ),
    .mux_select  ( set_muxes$029$mux_select ),
    .mux_out     ( set_muxes$029$mux_out )
  );

  // set_muxes$030 temporaries
  logic   [   5:0] set_muxes$030$mux_in_$000;
  logic   [   5:0] set_muxes$030$mux_in_$001;
  logic   [   0:0] set_muxes$030$clk;
  logic   [   0:0] set_muxes$030$reset;
  logic   [   0:0] set_muxes$030$mux_select;
  logic   [   5:0] set_muxes$030$mux_out;

  Mux_0x387678144da2c8e set_muxes$030
  (
    .mux_in_$000 ( set_muxes$030$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$030$mux_in_$001 ),
    .clk         ( set_muxes$030$clk ),
    .reset       ( set_muxes$030$reset ),
    .mux_select  ( set_muxes$030$mux_select ),
    .mux_out     ( set_muxes$030$mux_out )
  );

  // set_muxes$031 temporaries
  logic   [   5:0] set_muxes$031$mux_in_$000;
  logic   [   5:0] set_muxes$031$mux_in_$001;
  logic   [   0:0] set_muxes$031$clk;
  logic   [   0:0] set_muxes$031$reset;
  logic   [   0:0] set_muxes$031$mux_select;
  logic   [   5:0] set_muxes$031$mux_out;

  Mux_0x387678144da2c8e set_muxes$031
  (
    .mux_in_$000 ( set_muxes$031$mux_in_$000 ),
    .mux_in_$001 ( set_muxes$031$mux_in_$001 ),
    .clk         ( set_muxes$031$clk ),
    .reset       ( set_muxes$031$reset ),
    .mux_select  ( set_muxes$031$mux_select ),
    .mux_out     ( set_muxes$031$mux_out )
  );

  // snapshots$000 temporaries
  logic   [   5:0] snapshots$000$set_in_$000;
  logic   [   5:0] snapshots$000$set_in_$001;
  logic   [   5:0] snapshots$000$set_in_$002;
  logic   [   5:0] snapshots$000$set_in_$003;
  logic   [   5:0] snapshots$000$set_in_$004;
  logic   [   5:0] snapshots$000$set_in_$005;
  logic   [   5:0] snapshots$000$set_in_$006;
  logic   [   5:0] snapshots$000$set_in_$007;
  logic   [   5:0] snapshots$000$set_in_$008;
  logic   [   5:0] snapshots$000$set_in_$009;
  logic   [   5:0] snapshots$000$set_in_$010;
  logic   [   5:0] snapshots$000$set_in_$011;
  logic   [   5:0] snapshots$000$set_in_$012;
  logic   [   5:0] snapshots$000$set_in_$013;
  logic   [   5:0] snapshots$000$set_in_$014;
  logic   [   5:0] snapshots$000$set_in_$015;
  logic   [   5:0] snapshots$000$set_in_$016;
  logic   [   5:0] snapshots$000$set_in_$017;
  logic   [   5:0] snapshots$000$set_in_$018;
  logic   [   5:0] snapshots$000$set_in_$019;
  logic   [   5:0] snapshots$000$set_in_$020;
  logic   [   5:0] snapshots$000$set_in_$021;
  logic   [   5:0] snapshots$000$set_in_$022;
  logic   [   5:0] snapshots$000$set_in_$023;
  logic   [   5:0] snapshots$000$set_in_$024;
  logic   [   5:0] snapshots$000$set_in_$025;
  logic   [   5:0] snapshots$000$set_in_$026;
  logic   [   5:0] snapshots$000$set_in_$027;
  logic   [   5:0] snapshots$000$set_in_$028;
  logic   [   5:0] snapshots$000$set_in_$029;
  logic   [   5:0] snapshots$000$set_in_$030;
  logic   [   5:0] snapshots$000$set_in_$031;
  logic   [   0:0] snapshots$000$set_call;
  logic   [   0:0] snapshots$000$clk;
  logic   [   0:0] snapshots$000$reset;
  logic   [   5:0] snapshots$000$dump_out$000;
  logic   [   5:0] snapshots$000$dump_out$001;
  logic   [   5:0] snapshots$000$dump_out$002;
  logic   [   5:0] snapshots$000$dump_out$003;
  logic   [   5:0] snapshots$000$dump_out$004;
  logic   [   5:0] snapshots$000$dump_out$005;
  logic   [   5:0] snapshots$000$dump_out$006;
  logic   [   5:0] snapshots$000$dump_out$007;
  logic   [   5:0] snapshots$000$dump_out$008;
  logic   [   5:0] snapshots$000$dump_out$009;
  logic   [   5:0] snapshots$000$dump_out$010;
  logic   [   5:0] snapshots$000$dump_out$011;
  logic   [   5:0] snapshots$000$dump_out$012;
  logic   [   5:0] snapshots$000$dump_out$013;
  logic   [   5:0] snapshots$000$dump_out$014;
  logic   [   5:0] snapshots$000$dump_out$015;
  logic   [   5:0] snapshots$000$dump_out$016;
  logic   [   5:0] snapshots$000$dump_out$017;
  logic   [   5:0] snapshots$000$dump_out$018;
  logic   [   5:0] snapshots$000$dump_out$019;
  logic   [   5:0] snapshots$000$dump_out$020;
  logic   [   5:0] snapshots$000$dump_out$021;
  logic   [   5:0] snapshots$000$dump_out$022;
  logic   [   5:0] snapshots$000$dump_out$023;
  logic   [   5:0] snapshots$000$dump_out$024;
  logic   [   5:0] snapshots$000$dump_out$025;
  logic   [   5:0] snapshots$000$dump_out$026;
  logic   [   5:0] snapshots$000$dump_out$027;
  logic   [   5:0] snapshots$000$dump_out$028;
  logic   [   5:0] snapshots$000$dump_out$029;
  logic   [   5:0] snapshots$000$dump_out$030;
  logic   [   5:0] snapshots$000$dump_out$031;

  RegisterFile_0x5b973c72ce6092d snapshots$000
  (
    .set_in_$000  ( snapshots$000$set_in_$000 ),
    .set_in_$001  ( snapshots$000$set_in_$001 ),
    .set_in_$002  ( snapshots$000$set_in_$002 ),
    .set_in_$003  ( snapshots$000$set_in_$003 ),
    .set_in_$004  ( snapshots$000$set_in_$004 ),
    .set_in_$005  ( snapshots$000$set_in_$005 ),
    .set_in_$006  ( snapshots$000$set_in_$006 ),
    .set_in_$007  ( snapshots$000$set_in_$007 ),
    .set_in_$008  ( snapshots$000$set_in_$008 ),
    .set_in_$009  ( snapshots$000$set_in_$009 ),
    .set_in_$010  ( snapshots$000$set_in_$010 ),
    .set_in_$011  ( snapshots$000$set_in_$011 ),
    .set_in_$012  ( snapshots$000$set_in_$012 ),
    .set_in_$013  ( snapshots$000$set_in_$013 ),
    .set_in_$014  ( snapshots$000$set_in_$014 ),
    .set_in_$015  ( snapshots$000$set_in_$015 ),
    .set_in_$016  ( snapshots$000$set_in_$016 ),
    .set_in_$017  ( snapshots$000$set_in_$017 ),
    .set_in_$018  ( snapshots$000$set_in_$018 ),
    .set_in_$019  ( snapshots$000$set_in_$019 ),
    .set_in_$020  ( snapshots$000$set_in_$020 ),
    .set_in_$021  ( snapshots$000$set_in_$021 ),
    .set_in_$022  ( snapshots$000$set_in_$022 ),
    .set_in_$023  ( snapshots$000$set_in_$023 ),
    .set_in_$024  ( snapshots$000$set_in_$024 ),
    .set_in_$025  ( snapshots$000$set_in_$025 ),
    .set_in_$026  ( snapshots$000$set_in_$026 ),
    .set_in_$027  ( snapshots$000$set_in_$027 ),
    .set_in_$028  ( snapshots$000$set_in_$028 ),
    .set_in_$029  ( snapshots$000$set_in_$029 ),
    .set_in_$030  ( snapshots$000$set_in_$030 ),
    .set_in_$031  ( snapshots$000$set_in_$031 ),
    .set_call     ( snapshots$000$set_call ),
    .clk          ( snapshots$000$clk ),
    .reset        ( snapshots$000$reset ),
    .dump_out$000 ( snapshots$000$dump_out$000 ),
    .dump_out$001 ( snapshots$000$dump_out$001 ),
    .dump_out$002 ( snapshots$000$dump_out$002 ),
    .dump_out$003 ( snapshots$000$dump_out$003 ),
    .dump_out$004 ( snapshots$000$dump_out$004 ),
    .dump_out$005 ( snapshots$000$dump_out$005 ),
    .dump_out$006 ( snapshots$000$dump_out$006 ),
    .dump_out$007 ( snapshots$000$dump_out$007 ),
    .dump_out$008 ( snapshots$000$dump_out$008 ),
    .dump_out$009 ( snapshots$000$dump_out$009 ),
    .dump_out$010 ( snapshots$000$dump_out$010 ),
    .dump_out$011 ( snapshots$000$dump_out$011 ),
    .dump_out$012 ( snapshots$000$dump_out$012 ),
    .dump_out$013 ( snapshots$000$dump_out$013 ),
    .dump_out$014 ( snapshots$000$dump_out$014 ),
    .dump_out$015 ( snapshots$000$dump_out$015 ),
    .dump_out$016 ( snapshots$000$dump_out$016 ),
    .dump_out$017 ( snapshots$000$dump_out$017 ),
    .dump_out$018 ( snapshots$000$dump_out$018 ),
    .dump_out$019 ( snapshots$000$dump_out$019 ),
    .dump_out$020 ( snapshots$000$dump_out$020 ),
    .dump_out$021 ( snapshots$000$dump_out$021 ),
    .dump_out$022 ( snapshots$000$dump_out$022 ),
    .dump_out$023 ( snapshots$000$dump_out$023 ),
    .dump_out$024 ( snapshots$000$dump_out$024 ),
    .dump_out$025 ( snapshots$000$dump_out$025 ),
    .dump_out$026 ( snapshots$000$dump_out$026 ),
    .dump_out$027 ( snapshots$000$dump_out$027 ),
    .dump_out$028 ( snapshots$000$dump_out$028 ),
    .dump_out$029 ( snapshots$000$dump_out$029 ),
    .dump_out$030 ( snapshots$000$dump_out$030 ),
    .dump_out$031 ( snapshots$000$dump_out$031 )
  );

  // snapshots$001 temporaries
  logic   [   5:0] snapshots$001$set_in_$000;
  logic   [   5:0] snapshots$001$set_in_$001;
  logic   [   5:0] snapshots$001$set_in_$002;
  logic   [   5:0] snapshots$001$set_in_$003;
  logic   [   5:0] snapshots$001$set_in_$004;
  logic   [   5:0] snapshots$001$set_in_$005;
  logic   [   5:0] snapshots$001$set_in_$006;
  logic   [   5:0] snapshots$001$set_in_$007;
  logic   [   5:0] snapshots$001$set_in_$008;
  logic   [   5:0] snapshots$001$set_in_$009;
  logic   [   5:0] snapshots$001$set_in_$010;
  logic   [   5:0] snapshots$001$set_in_$011;
  logic   [   5:0] snapshots$001$set_in_$012;
  logic   [   5:0] snapshots$001$set_in_$013;
  logic   [   5:0] snapshots$001$set_in_$014;
  logic   [   5:0] snapshots$001$set_in_$015;
  logic   [   5:0] snapshots$001$set_in_$016;
  logic   [   5:0] snapshots$001$set_in_$017;
  logic   [   5:0] snapshots$001$set_in_$018;
  logic   [   5:0] snapshots$001$set_in_$019;
  logic   [   5:0] snapshots$001$set_in_$020;
  logic   [   5:0] snapshots$001$set_in_$021;
  logic   [   5:0] snapshots$001$set_in_$022;
  logic   [   5:0] snapshots$001$set_in_$023;
  logic   [   5:0] snapshots$001$set_in_$024;
  logic   [   5:0] snapshots$001$set_in_$025;
  logic   [   5:0] snapshots$001$set_in_$026;
  logic   [   5:0] snapshots$001$set_in_$027;
  logic   [   5:0] snapshots$001$set_in_$028;
  logic   [   5:0] snapshots$001$set_in_$029;
  logic   [   5:0] snapshots$001$set_in_$030;
  logic   [   5:0] snapshots$001$set_in_$031;
  logic   [   0:0] snapshots$001$set_call;
  logic   [   0:0] snapshots$001$clk;
  logic   [   0:0] snapshots$001$reset;
  logic   [   5:0] snapshots$001$dump_out$000;
  logic   [   5:0] snapshots$001$dump_out$001;
  logic   [   5:0] snapshots$001$dump_out$002;
  logic   [   5:0] snapshots$001$dump_out$003;
  logic   [   5:0] snapshots$001$dump_out$004;
  logic   [   5:0] snapshots$001$dump_out$005;
  logic   [   5:0] snapshots$001$dump_out$006;
  logic   [   5:0] snapshots$001$dump_out$007;
  logic   [   5:0] snapshots$001$dump_out$008;
  logic   [   5:0] snapshots$001$dump_out$009;
  logic   [   5:0] snapshots$001$dump_out$010;
  logic   [   5:0] snapshots$001$dump_out$011;
  logic   [   5:0] snapshots$001$dump_out$012;
  logic   [   5:0] snapshots$001$dump_out$013;
  logic   [   5:0] snapshots$001$dump_out$014;
  logic   [   5:0] snapshots$001$dump_out$015;
  logic   [   5:0] snapshots$001$dump_out$016;
  logic   [   5:0] snapshots$001$dump_out$017;
  logic   [   5:0] snapshots$001$dump_out$018;
  logic   [   5:0] snapshots$001$dump_out$019;
  logic   [   5:0] snapshots$001$dump_out$020;
  logic   [   5:0] snapshots$001$dump_out$021;
  logic   [   5:0] snapshots$001$dump_out$022;
  logic   [   5:0] snapshots$001$dump_out$023;
  logic   [   5:0] snapshots$001$dump_out$024;
  logic   [   5:0] snapshots$001$dump_out$025;
  logic   [   5:0] snapshots$001$dump_out$026;
  logic   [   5:0] snapshots$001$dump_out$027;
  logic   [   5:0] snapshots$001$dump_out$028;
  logic   [   5:0] snapshots$001$dump_out$029;
  logic   [   5:0] snapshots$001$dump_out$030;
  logic   [   5:0] snapshots$001$dump_out$031;

  RegisterFile_0x5b973c72ce6092d snapshots$001
  (
    .set_in_$000  ( snapshots$001$set_in_$000 ),
    .set_in_$001  ( snapshots$001$set_in_$001 ),
    .set_in_$002  ( snapshots$001$set_in_$002 ),
    .set_in_$003  ( snapshots$001$set_in_$003 ),
    .set_in_$004  ( snapshots$001$set_in_$004 ),
    .set_in_$005  ( snapshots$001$set_in_$005 ),
    .set_in_$006  ( snapshots$001$set_in_$006 ),
    .set_in_$007  ( snapshots$001$set_in_$007 ),
    .set_in_$008  ( snapshots$001$set_in_$008 ),
    .set_in_$009  ( snapshots$001$set_in_$009 ),
    .set_in_$010  ( snapshots$001$set_in_$010 ),
    .set_in_$011  ( snapshots$001$set_in_$011 ),
    .set_in_$012  ( snapshots$001$set_in_$012 ),
    .set_in_$013  ( snapshots$001$set_in_$013 ),
    .set_in_$014  ( snapshots$001$set_in_$014 ),
    .set_in_$015  ( snapshots$001$set_in_$015 ),
    .set_in_$016  ( snapshots$001$set_in_$016 ),
    .set_in_$017  ( snapshots$001$set_in_$017 ),
    .set_in_$018  ( snapshots$001$set_in_$018 ),
    .set_in_$019  ( snapshots$001$set_in_$019 ),
    .set_in_$020  ( snapshots$001$set_in_$020 ),
    .set_in_$021  ( snapshots$001$set_in_$021 ),
    .set_in_$022  ( snapshots$001$set_in_$022 ),
    .set_in_$023  ( snapshots$001$set_in_$023 ),
    .set_in_$024  ( snapshots$001$set_in_$024 ),
    .set_in_$025  ( snapshots$001$set_in_$025 ),
    .set_in_$026  ( snapshots$001$set_in_$026 ),
    .set_in_$027  ( snapshots$001$set_in_$027 ),
    .set_in_$028  ( snapshots$001$set_in_$028 ),
    .set_in_$029  ( snapshots$001$set_in_$029 ),
    .set_in_$030  ( snapshots$001$set_in_$030 ),
    .set_in_$031  ( snapshots$001$set_in_$031 ),
    .set_call     ( snapshots$001$set_call ),
    .clk          ( snapshots$001$clk ),
    .reset        ( snapshots$001$reset ),
    .dump_out$000 ( snapshots$001$dump_out$000 ),
    .dump_out$001 ( snapshots$001$dump_out$001 ),
    .dump_out$002 ( snapshots$001$dump_out$002 ),
    .dump_out$003 ( snapshots$001$dump_out$003 ),
    .dump_out$004 ( snapshots$001$dump_out$004 ),
    .dump_out$005 ( snapshots$001$dump_out$005 ),
    .dump_out$006 ( snapshots$001$dump_out$006 ),
    .dump_out$007 ( snapshots$001$dump_out$007 ),
    .dump_out$008 ( snapshots$001$dump_out$008 ),
    .dump_out$009 ( snapshots$001$dump_out$009 ),
    .dump_out$010 ( snapshots$001$dump_out$010 ),
    .dump_out$011 ( snapshots$001$dump_out$011 ),
    .dump_out$012 ( snapshots$001$dump_out$012 ),
    .dump_out$013 ( snapshots$001$dump_out$013 ),
    .dump_out$014 ( snapshots$001$dump_out$014 ),
    .dump_out$015 ( snapshots$001$dump_out$015 ),
    .dump_out$016 ( snapshots$001$dump_out$016 ),
    .dump_out$017 ( snapshots$001$dump_out$017 ),
    .dump_out$018 ( snapshots$001$dump_out$018 ),
    .dump_out$019 ( snapshots$001$dump_out$019 ),
    .dump_out$020 ( snapshots$001$dump_out$020 ),
    .dump_out$021 ( snapshots$001$dump_out$021 ),
    .dump_out$022 ( snapshots$001$dump_out$022 ),
    .dump_out$023 ( snapshots$001$dump_out$023 ),
    .dump_out$024 ( snapshots$001$dump_out$024 ),
    .dump_out$025 ( snapshots$001$dump_out$025 ),
    .dump_out$026 ( snapshots$001$dump_out$026 ),
    .dump_out$027 ( snapshots$001$dump_out$027 ),
    .dump_out$028 ( snapshots$001$dump_out$028 ),
    .dump_out$029 ( snapshots$001$dump_out$029 ),
    .dump_out$030 ( snapshots$001$dump_out$030 ),
    .dump_out$031 ( snapshots$001$dump_out$031 )
  );

  // signal connections
  assign read_data$000                  = regs$read_data$000;
  assign read_data$001                  = regs$read_data$001;
  assign regs$clk                       = clk;
  assign regs$read_addr$000             = read_addr$000;
  assign regs$read_addr$001             = read_addr$001;
  assign regs$reset                     = reset;
  assign regs$set_call                  = should_set;
  assign regs$set_in_$000               = set_muxes$000$mux_out;
  assign regs$set_in_$001               = set_muxes$001$mux_out;
  assign regs$set_in_$002               = set_muxes$002$mux_out;
  assign regs$set_in_$003               = set_muxes$003$mux_out;
  assign regs$set_in_$004               = set_muxes$004$mux_out;
  assign regs$set_in_$005               = set_muxes$005$mux_out;
  assign regs$set_in_$006               = set_muxes$006$mux_out;
  assign regs$set_in_$007               = set_muxes$007$mux_out;
  assign regs$set_in_$008               = set_muxes$008$mux_out;
  assign regs$set_in_$009               = set_muxes$009$mux_out;
  assign regs$set_in_$010               = set_muxes$010$mux_out;
  assign regs$set_in_$011               = set_muxes$011$mux_out;
  assign regs$set_in_$012               = set_muxes$012$mux_out;
  assign regs$set_in_$013               = set_muxes$013$mux_out;
  assign regs$set_in_$014               = set_muxes$014$mux_out;
  assign regs$set_in_$015               = set_muxes$015$mux_out;
  assign regs$set_in_$016               = set_muxes$016$mux_out;
  assign regs$set_in_$017               = set_muxes$017$mux_out;
  assign regs$set_in_$018               = set_muxes$018$mux_out;
  assign regs$set_in_$019               = set_muxes$019$mux_out;
  assign regs$set_in_$020               = set_muxes$020$mux_out;
  assign regs$set_in_$021               = set_muxes$021$mux_out;
  assign regs$set_in_$022               = set_muxes$022$mux_out;
  assign regs$set_in_$023               = set_muxes$023$mux_out;
  assign regs$set_in_$024               = set_muxes$024$mux_out;
  assign regs$set_in_$025               = set_muxes$025$mux_out;
  assign regs$set_in_$026               = set_muxes$026$mux_out;
  assign regs$set_in_$027               = set_muxes$027$mux_out;
  assign regs$set_in_$028               = set_muxes$028$mux_out;
  assign regs$set_in_$029               = set_muxes$029$mux_out;
  assign regs$set_in_$030               = set_muxes$030$mux_out;
  assign regs$set_in_$031               = set_muxes$031$mux_out;
  assign regs$write_addr$000            = write_addr$000;
  assign regs$write_call$000            = write_call$000;
  assign regs$write_data$000            = write_data$000;
  assign restore_vector$000             = snapshot_muxes$000$mux_out;
  assign restore_vector$001             = snapshot_muxes$001$mux_out;
  assign restore_vector$002             = snapshot_muxes$002$mux_out;
  assign restore_vector$003             = snapshot_muxes$003$mux_out;
  assign restore_vector$004             = snapshot_muxes$004$mux_out;
  assign restore_vector$005             = snapshot_muxes$005$mux_out;
  assign restore_vector$006             = snapshot_muxes$006$mux_out;
  assign restore_vector$007             = snapshot_muxes$007$mux_out;
  assign restore_vector$008             = snapshot_muxes$008$mux_out;
  assign restore_vector$009             = snapshot_muxes$009$mux_out;
  assign restore_vector$010             = snapshot_muxes$010$mux_out;
  assign restore_vector$011             = snapshot_muxes$011$mux_out;
  assign restore_vector$012             = snapshot_muxes$012$mux_out;
  assign restore_vector$013             = snapshot_muxes$013$mux_out;
  assign restore_vector$014             = snapshot_muxes$014$mux_out;
  assign restore_vector$015             = snapshot_muxes$015$mux_out;
  assign restore_vector$016             = snapshot_muxes$016$mux_out;
  assign restore_vector$017             = snapshot_muxes$017$mux_out;
  assign restore_vector$018             = snapshot_muxes$018$mux_out;
  assign restore_vector$019             = snapshot_muxes$019$mux_out;
  assign restore_vector$020             = snapshot_muxes$020$mux_out;
  assign restore_vector$021             = snapshot_muxes$021$mux_out;
  assign restore_vector$022             = snapshot_muxes$022$mux_out;
  assign restore_vector$023             = snapshot_muxes$023$mux_out;
  assign restore_vector$024             = snapshot_muxes$024$mux_out;
  assign restore_vector$025             = snapshot_muxes$025$mux_out;
  assign restore_vector$026             = snapshot_muxes$026$mux_out;
  assign restore_vector$027             = snapshot_muxes$027$mux_out;
  assign restore_vector$028             = snapshot_muxes$028$mux_out;
  assign restore_vector$029             = snapshot_muxes$029$mux_out;
  assign restore_vector$030             = snapshot_muxes$030$mux_out;
  assign restore_vector$031             = snapshot_muxes$031$mux_out;
  assign set_muxes$000$clk              = clk;
  assign set_muxes$000$mux_in_$000      = restore_vector$000;
  assign set_muxes$000$mux_in_$001      = set_in_$000;
  assign set_muxes$000$mux_select       = set_call;
  assign set_muxes$000$reset            = reset;
  assign set_muxes$001$clk              = clk;
  assign set_muxes$001$mux_in_$000      = restore_vector$001;
  assign set_muxes$001$mux_in_$001      = set_in_$001;
  assign set_muxes$001$mux_select       = set_call;
  assign set_muxes$001$reset            = reset;
  assign set_muxes$002$clk              = clk;
  assign set_muxes$002$mux_in_$000      = restore_vector$002;
  assign set_muxes$002$mux_in_$001      = set_in_$002;
  assign set_muxes$002$mux_select       = set_call;
  assign set_muxes$002$reset            = reset;
  assign set_muxes$003$clk              = clk;
  assign set_muxes$003$mux_in_$000      = restore_vector$003;
  assign set_muxes$003$mux_in_$001      = set_in_$003;
  assign set_muxes$003$mux_select       = set_call;
  assign set_muxes$003$reset            = reset;
  assign set_muxes$004$clk              = clk;
  assign set_muxes$004$mux_in_$000      = restore_vector$004;
  assign set_muxes$004$mux_in_$001      = set_in_$004;
  assign set_muxes$004$mux_select       = set_call;
  assign set_muxes$004$reset            = reset;
  assign set_muxes$005$clk              = clk;
  assign set_muxes$005$mux_in_$000      = restore_vector$005;
  assign set_muxes$005$mux_in_$001      = set_in_$005;
  assign set_muxes$005$mux_select       = set_call;
  assign set_muxes$005$reset            = reset;
  assign set_muxes$006$clk              = clk;
  assign set_muxes$006$mux_in_$000      = restore_vector$006;
  assign set_muxes$006$mux_in_$001      = set_in_$006;
  assign set_muxes$006$mux_select       = set_call;
  assign set_muxes$006$reset            = reset;
  assign set_muxes$007$clk              = clk;
  assign set_muxes$007$mux_in_$000      = restore_vector$007;
  assign set_muxes$007$mux_in_$001      = set_in_$007;
  assign set_muxes$007$mux_select       = set_call;
  assign set_muxes$007$reset            = reset;
  assign set_muxes$008$clk              = clk;
  assign set_muxes$008$mux_in_$000      = restore_vector$008;
  assign set_muxes$008$mux_in_$001      = set_in_$008;
  assign set_muxes$008$mux_select       = set_call;
  assign set_muxes$008$reset            = reset;
  assign set_muxes$009$clk              = clk;
  assign set_muxes$009$mux_in_$000      = restore_vector$009;
  assign set_muxes$009$mux_in_$001      = set_in_$009;
  assign set_muxes$009$mux_select       = set_call;
  assign set_muxes$009$reset            = reset;
  assign set_muxes$010$clk              = clk;
  assign set_muxes$010$mux_in_$000      = restore_vector$010;
  assign set_muxes$010$mux_in_$001      = set_in_$010;
  assign set_muxes$010$mux_select       = set_call;
  assign set_muxes$010$reset            = reset;
  assign set_muxes$011$clk              = clk;
  assign set_muxes$011$mux_in_$000      = restore_vector$011;
  assign set_muxes$011$mux_in_$001      = set_in_$011;
  assign set_muxes$011$mux_select       = set_call;
  assign set_muxes$011$reset            = reset;
  assign set_muxes$012$clk              = clk;
  assign set_muxes$012$mux_in_$000      = restore_vector$012;
  assign set_muxes$012$mux_in_$001      = set_in_$012;
  assign set_muxes$012$mux_select       = set_call;
  assign set_muxes$012$reset            = reset;
  assign set_muxes$013$clk              = clk;
  assign set_muxes$013$mux_in_$000      = restore_vector$013;
  assign set_muxes$013$mux_in_$001      = set_in_$013;
  assign set_muxes$013$mux_select       = set_call;
  assign set_muxes$013$reset            = reset;
  assign set_muxes$014$clk              = clk;
  assign set_muxes$014$mux_in_$000      = restore_vector$014;
  assign set_muxes$014$mux_in_$001      = set_in_$014;
  assign set_muxes$014$mux_select       = set_call;
  assign set_muxes$014$reset            = reset;
  assign set_muxes$015$clk              = clk;
  assign set_muxes$015$mux_in_$000      = restore_vector$015;
  assign set_muxes$015$mux_in_$001      = set_in_$015;
  assign set_muxes$015$mux_select       = set_call;
  assign set_muxes$015$reset            = reset;
  assign set_muxes$016$clk              = clk;
  assign set_muxes$016$mux_in_$000      = restore_vector$016;
  assign set_muxes$016$mux_in_$001      = set_in_$016;
  assign set_muxes$016$mux_select       = set_call;
  assign set_muxes$016$reset            = reset;
  assign set_muxes$017$clk              = clk;
  assign set_muxes$017$mux_in_$000      = restore_vector$017;
  assign set_muxes$017$mux_in_$001      = set_in_$017;
  assign set_muxes$017$mux_select       = set_call;
  assign set_muxes$017$reset            = reset;
  assign set_muxes$018$clk              = clk;
  assign set_muxes$018$mux_in_$000      = restore_vector$018;
  assign set_muxes$018$mux_in_$001      = set_in_$018;
  assign set_muxes$018$mux_select       = set_call;
  assign set_muxes$018$reset            = reset;
  assign set_muxes$019$clk              = clk;
  assign set_muxes$019$mux_in_$000      = restore_vector$019;
  assign set_muxes$019$mux_in_$001      = set_in_$019;
  assign set_muxes$019$mux_select       = set_call;
  assign set_muxes$019$reset            = reset;
  assign set_muxes$020$clk              = clk;
  assign set_muxes$020$mux_in_$000      = restore_vector$020;
  assign set_muxes$020$mux_in_$001      = set_in_$020;
  assign set_muxes$020$mux_select       = set_call;
  assign set_muxes$020$reset            = reset;
  assign set_muxes$021$clk              = clk;
  assign set_muxes$021$mux_in_$000      = restore_vector$021;
  assign set_muxes$021$mux_in_$001      = set_in_$021;
  assign set_muxes$021$mux_select       = set_call;
  assign set_muxes$021$reset            = reset;
  assign set_muxes$022$clk              = clk;
  assign set_muxes$022$mux_in_$000      = restore_vector$022;
  assign set_muxes$022$mux_in_$001      = set_in_$022;
  assign set_muxes$022$mux_select       = set_call;
  assign set_muxes$022$reset            = reset;
  assign set_muxes$023$clk              = clk;
  assign set_muxes$023$mux_in_$000      = restore_vector$023;
  assign set_muxes$023$mux_in_$001      = set_in_$023;
  assign set_muxes$023$mux_select       = set_call;
  assign set_muxes$023$reset            = reset;
  assign set_muxes$024$clk              = clk;
  assign set_muxes$024$mux_in_$000      = restore_vector$024;
  assign set_muxes$024$mux_in_$001      = set_in_$024;
  assign set_muxes$024$mux_select       = set_call;
  assign set_muxes$024$reset            = reset;
  assign set_muxes$025$clk              = clk;
  assign set_muxes$025$mux_in_$000      = restore_vector$025;
  assign set_muxes$025$mux_in_$001      = set_in_$025;
  assign set_muxes$025$mux_select       = set_call;
  assign set_muxes$025$reset            = reset;
  assign set_muxes$026$clk              = clk;
  assign set_muxes$026$mux_in_$000      = restore_vector$026;
  assign set_muxes$026$mux_in_$001      = set_in_$026;
  assign set_muxes$026$mux_select       = set_call;
  assign set_muxes$026$reset            = reset;
  assign set_muxes$027$clk              = clk;
  assign set_muxes$027$mux_in_$000      = restore_vector$027;
  assign set_muxes$027$mux_in_$001      = set_in_$027;
  assign set_muxes$027$mux_select       = set_call;
  assign set_muxes$027$reset            = reset;
  assign set_muxes$028$clk              = clk;
  assign set_muxes$028$mux_in_$000      = restore_vector$028;
  assign set_muxes$028$mux_in_$001      = set_in_$028;
  assign set_muxes$028$mux_select       = set_call;
  assign set_muxes$028$reset            = reset;
  assign set_muxes$029$clk              = clk;
  assign set_muxes$029$mux_in_$000      = restore_vector$029;
  assign set_muxes$029$mux_in_$001      = set_in_$029;
  assign set_muxes$029$mux_select       = set_call;
  assign set_muxes$029$reset            = reset;
  assign set_muxes$030$clk              = clk;
  assign set_muxes$030$mux_in_$000      = restore_vector$030;
  assign set_muxes$030$mux_in_$001      = set_in_$030;
  assign set_muxes$030$mux_select       = set_call;
  assign set_muxes$030$reset            = reset;
  assign set_muxes$031$clk              = clk;
  assign set_muxes$031$mux_in_$000      = restore_vector$031;
  assign set_muxes$031$mux_in_$001      = set_in_$031;
  assign set_muxes$031$mux_select       = set_call;
  assign set_muxes$031$reset            = reset;
  assign snapshot_muxes$000$clk         = clk;
  assign snapshot_muxes$000$mux_in_$000 = snapshots$000$dump_out$000;
  assign snapshot_muxes$000$mux_in_$001 = snapshots$001$dump_out$000;
  assign snapshot_muxes$000$mux_select  = restore_source_id;
  assign snapshot_muxes$000$reset       = reset;
  assign snapshot_muxes$001$clk         = clk;
  assign snapshot_muxes$001$mux_in_$000 = snapshots$000$dump_out$001;
  assign snapshot_muxes$001$mux_in_$001 = snapshots$001$dump_out$001;
  assign snapshot_muxes$001$mux_select  = restore_source_id;
  assign snapshot_muxes$001$reset       = reset;
  assign snapshot_muxes$002$clk         = clk;
  assign snapshot_muxes$002$mux_in_$000 = snapshots$000$dump_out$002;
  assign snapshot_muxes$002$mux_in_$001 = snapshots$001$dump_out$002;
  assign snapshot_muxes$002$mux_select  = restore_source_id;
  assign snapshot_muxes$002$reset       = reset;
  assign snapshot_muxes$003$clk         = clk;
  assign snapshot_muxes$003$mux_in_$000 = snapshots$000$dump_out$003;
  assign snapshot_muxes$003$mux_in_$001 = snapshots$001$dump_out$003;
  assign snapshot_muxes$003$mux_select  = restore_source_id;
  assign snapshot_muxes$003$reset       = reset;
  assign snapshot_muxes$004$clk         = clk;
  assign snapshot_muxes$004$mux_in_$000 = snapshots$000$dump_out$004;
  assign snapshot_muxes$004$mux_in_$001 = snapshots$001$dump_out$004;
  assign snapshot_muxes$004$mux_select  = restore_source_id;
  assign snapshot_muxes$004$reset       = reset;
  assign snapshot_muxes$005$clk         = clk;
  assign snapshot_muxes$005$mux_in_$000 = snapshots$000$dump_out$005;
  assign snapshot_muxes$005$mux_in_$001 = snapshots$001$dump_out$005;
  assign snapshot_muxes$005$mux_select  = restore_source_id;
  assign snapshot_muxes$005$reset       = reset;
  assign snapshot_muxes$006$clk         = clk;
  assign snapshot_muxes$006$mux_in_$000 = snapshots$000$dump_out$006;
  assign snapshot_muxes$006$mux_in_$001 = snapshots$001$dump_out$006;
  assign snapshot_muxes$006$mux_select  = restore_source_id;
  assign snapshot_muxes$006$reset       = reset;
  assign snapshot_muxes$007$clk         = clk;
  assign snapshot_muxes$007$mux_in_$000 = snapshots$000$dump_out$007;
  assign snapshot_muxes$007$mux_in_$001 = snapshots$001$dump_out$007;
  assign snapshot_muxes$007$mux_select  = restore_source_id;
  assign snapshot_muxes$007$reset       = reset;
  assign snapshot_muxes$008$clk         = clk;
  assign snapshot_muxes$008$mux_in_$000 = snapshots$000$dump_out$008;
  assign snapshot_muxes$008$mux_in_$001 = snapshots$001$dump_out$008;
  assign snapshot_muxes$008$mux_select  = restore_source_id;
  assign snapshot_muxes$008$reset       = reset;
  assign snapshot_muxes$009$clk         = clk;
  assign snapshot_muxes$009$mux_in_$000 = snapshots$000$dump_out$009;
  assign snapshot_muxes$009$mux_in_$001 = snapshots$001$dump_out$009;
  assign snapshot_muxes$009$mux_select  = restore_source_id;
  assign snapshot_muxes$009$reset       = reset;
  assign snapshot_muxes$010$clk         = clk;
  assign snapshot_muxes$010$mux_in_$000 = snapshots$000$dump_out$010;
  assign snapshot_muxes$010$mux_in_$001 = snapshots$001$dump_out$010;
  assign snapshot_muxes$010$mux_select  = restore_source_id;
  assign snapshot_muxes$010$reset       = reset;
  assign snapshot_muxes$011$clk         = clk;
  assign snapshot_muxes$011$mux_in_$000 = snapshots$000$dump_out$011;
  assign snapshot_muxes$011$mux_in_$001 = snapshots$001$dump_out$011;
  assign snapshot_muxes$011$mux_select  = restore_source_id;
  assign snapshot_muxes$011$reset       = reset;
  assign snapshot_muxes$012$clk         = clk;
  assign snapshot_muxes$012$mux_in_$000 = snapshots$000$dump_out$012;
  assign snapshot_muxes$012$mux_in_$001 = snapshots$001$dump_out$012;
  assign snapshot_muxes$012$mux_select  = restore_source_id;
  assign snapshot_muxes$012$reset       = reset;
  assign snapshot_muxes$013$clk         = clk;
  assign snapshot_muxes$013$mux_in_$000 = snapshots$000$dump_out$013;
  assign snapshot_muxes$013$mux_in_$001 = snapshots$001$dump_out$013;
  assign snapshot_muxes$013$mux_select  = restore_source_id;
  assign snapshot_muxes$013$reset       = reset;
  assign snapshot_muxes$014$clk         = clk;
  assign snapshot_muxes$014$mux_in_$000 = snapshots$000$dump_out$014;
  assign snapshot_muxes$014$mux_in_$001 = snapshots$001$dump_out$014;
  assign snapshot_muxes$014$mux_select  = restore_source_id;
  assign snapshot_muxes$014$reset       = reset;
  assign snapshot_muxes$015$clk         = clk;
  assign snapshot_muxes$015$mux_in_$000 = snapshots$000$dump_out$015;
  assign snapshot_muxes$015$mux_in_$001 = snapshots$001$dump_out$015;
  assign snapshot_muxes$015$mux_select  = restore_source_id;
  assign snapshot_muxes$015$reset       = reset;
  assign snapshot_muxes$016$clk         = clk;
  assign snapshot_muxes$016$mux_in_$000 = snapshots$000$dump_out$016;
  assign snapshot_muxes$016$mux_in_$001 = snapshots$001$dump_out$016;
  assign snapshot_muxes$016$mux_select  = restore_source_id;
  assign snapshot_muxes$016$reset       = reset;
  assign snapshot_muxes$017$clk         = clk;
  assign snapshot_muxes$017$mux_in_$000 = snapshots$000$dump_out$017;
  assign snapshot_muxes$017$mux_in_$001 = snapshots$001$dump_out$017;
  assign snapshot_muxes$017$mux_select  = restore_source_id;
  assign snapshot_muxes$017$reset       = reset;
  assign snapshot_muxes$018$clk         = clk;
  assign snapshot_muxes$018$mux_in_$000 = snapshots$000$dump_out$018;
  assign snapshot_muxes$018$mux_in_$001 = snapshots$001$dump_out$018;
  assign snapshot_muxes$018$mux_select  = restore_source_id;
  assign snapshot_muxes$018$reset       = reset;
  assign snapshot_muxes$019$clk         = clk;
  assign snapshot_muxes$019$mux_in_$000 = snapshots$000$dump_out$019;
  assign snapshot_muxes$019$mux_in_$001 = snapshots$001$dump_out$019;
  assign snapshot_muxes$019$mux_select  = restore_source_id;
  assign snapshot_muxes$019$reset       = reset;
  assign snapshot_muxes$020$clk         = clk;
  assign snapshot_muxes$020$mux_in_$000 = snapshots$000$dump_out$020;
  assign snapshot_muxes$020$mux_in_$001 = snapshots$001$dump_out$020;
  assign snapshot_muxes$020$mux_select  = restore_source_id;
  assign snapshot_muxes$020$reset       = reset;
  assign snapshot_muxes$021$clk         = clk;
  assign snapshot_muxes$021$mux_in_$000 = snapshots$000$dump_out$021;
  assign snapshot_muxes$021$mux_in_$001 = snapshots$001$dump_out$021;
  assign snapshot_muxes$021$mux_select  = restore_source_id;
  assign snapshot_muxes$021$reset       = reset;
  assign snapshot_muxes$022$clk         = clk;
  assign snapshot_muxes$022$mux_in_$000 = snapshots$000$dump_out$022;
  assign snapshot_muxes$022$mux_in_$001 = snapshots$001$dump_out$022;
  assign snapshot_muxes$022$mux_select  = restore_source_id;
  assign snapshot_muxes$022$reset       = reset;
  assign snapshot_muxes$023$clk         = clk;
  assign snapshot_muxes$023$mux_in_$000 = snapshots$000$dump_out$023;
  assign snapshot_muxes$023$mux_in_$001 = snapshots$001$dump_out$023;
  assign snapshot_muxes$023$mux_select  = restore_source_id;
  assign snapshot_muxes$023$reset       = reset;
  assign snapshot_muxes$024$clk         = clk;
  assign snapshot_muxes$024$mux_in_$000 = snapshots$000$dump_out$024;
  assign snapshot_muxes$024$mux_in_$001 = snapshots$001$dump_out$024;
  assign snapshot_muxes$024$mux_select  = restore_source_id;
  assign snapshot_muxes$024$reset       = reset;
  assign snapshot_muxes$025$clk         = clk;
  assign snapshot_muxes$025$mux_in_$000 = snapshots$000$dump_out$025;
  assign snapshot_muxes$025$mux_in_$001 = snapshots$001$dump_out$025;
  assign snapshot_muxes$025$mux_select  = restore_source_id;
  assign snapshot_muxes$025$reset       = reset;
  assign snapshot_muxes$026$clk         = clk;
  assign snapshot_muxes$026$mux_in_$000 = snapshots$000$dump_out$026;
  assign snapshot_muxes$026$mux_in_$001 = snapshots$001$dump_out$026;
  assign snapshot_muxes$026$mux_select  = restore_source_id;
  assign snapshot_muxes$026$reset       = reset;
  assign snapshot_muxes$027$clk         = clk;
  assign snapshot_muxes$027$mux_in_$000 = snapshots$000$dump_out$027;
  assign snapshot_muxes$027$mux_in_$001 = snapshots$001$dump_out$027;
  assign snapshot_muxes$027$mux_select  = restore_source_id;
  assign snapshot_muxes$027$reset       = reset;
  assign snapshot_muxes$028$clk         = clk;
  assign snapshot_muxes$028$mux_in_$000 = snapshots$000$dump_out$028;
  assign snapshot_muxes$028$mux_in_$001 = snapshots$001$dump_out$028;
  assign snapshot_muxes$028$mux_select  = restore_source_id;
  assign snapshot_muxes$028$reset       = reset;
  assign snapshot_muxes$029$clk         = clk;
  assign snapshot_muxes$029$mux_in_$000 = snapshots$000$dump_out$029;
  assign snapshot_muxes$029$mux_in_$001 = snapshots$001$dump_out$029;
  assign snapshot_muxes$029$mux_select  = restore_source_id;
  assign snapshot_muxes$029$reset       = reset;
  assign snapshot_muxes$030$clk         = clk;
  assign snapshot_muxes$030$mux_in_$000 = snapshots$000$dump_out$030;
  assign snapshot_muxes$030$mux_in_$001 = snapshots$001$dump_out$030;
  assign snapshot_muxes$030$mux_select  = restore_source_id;
  assign snapshot_muxes$030$reset       = reset;
  assign snapshot_muxes$031$clk         = clk;
  assign snapshot_muxes$031$mux_in_$000 = snapshots$000$dump_out$031;
  assign snapshot_muxes$031$mux_in_$001 = snapshots$001$dump_out$031;
  assign snapshot_muxes$031$mux_select  = restore_source_id;
  assign snapshot_muxes$031$reset       = reset;
  assign snapshots$000$clk              = clk;
  assign snapshots$000$reset            = reset;
  assign snapshots$000$set_in_$000      = regs$dump_out$000;
  assign snapshots$000$set_in_$001      = regs$dump_out$001;
  assign snapshots$000$set_in_$002      = regs$dump_out$002;
  assign snapshots$000$set_in_$003      = regs$dump_out$003;
  assign snapshots$000$set_in_$004      = regs$dump_out$004;
  assign snapshots$000$set_in_$005      = regs$dump_out$005;
  assign snapshots$000$set_in_$006      = regs$dump_out$006;
  assign snapshots$000$set_in_$007      = regs$dump_out$007;
  assign snapshots$000$set_in_$008      = regs$dump_out$008;
  assign snapshots$000$set_in_$009      = regs$dump_out$009;
  assign snapshots$000$set_in_$010      = regs$dump_out$010;
  assign snapshots$000$set_in_$011      = regs$dump_out$011;
  assign snapshots$000$set_in_$012      = regs$dump_out$012;
  assign snapshots$000$set_in_$013      = regs$dump_out$013;
  assign snapshots$000$set_in_$014      = regs$dump_out$014;
  assign snapshots$000$set_in_$015      = regs$dump_out$015;
  assign snapshots$000$set_in_$016      = regs$dump_out$016;
  assign snapshots$000$set_in_$017      = regs$dump_out$017;
  assign snapshots$000$set_in_$018      = regs$dump_out$018;
  assign snapshots$000$set_in_$019      = regs$dump_out$019;
  assign snapshots$000$set_in_$020      = regs$dump_out$020;
  assign snapshots$000$set_in_$021      = regs$dump_out$021;
  assign snapshots$000$set_in_$022      = regs$dump_out$022;
  assign snapshots$000$set_in_$023      = regs$dump_out$023;
  assign snapshots$000$set_in_$024      = regs$dump_out$024;
  assign snapshots$000$set_in_$025      = regs$dump_out$025;
  assign snapshots$000$set_in_$026      = regs$dump_out$026;
  assign snapshots$000$set_in_$027      = regs$dump_out$027;
  assign snapshots$000$set_in_$028      = regs$dump_out$028;
  assign snapshots$000$set_in_$029      = regs$dump_out$029;
  assign snapshots$000$set_in_$030      = regs$dump_out$030;
  assign snapshots$000$set_in_$031      = regs$dump_out$031;
  assign snapshots$001$clk              = clk;
  assign snapshots$001$reset            = reset;
  assign snapshots$001$set_in_$000      = regs$dump_out$000;
  assign snapshots$001$set_in_$001      = regs$dump_out$001;
  assign snapshots$001$set_in_$002      = regs$dump_out$002;
  assign snapshots$001$set_in_$003      = regs$dump_out$003;
  assign snapshots$001$set_in_$004      = regs$dump_out$004;
  assign snapshots$001$set_in_$005      = regs$dump_out$005;
  assign snapshots$001$set_in_$006      = regs$dump_out$006;
  assign snapshots$001$set_in_$007      = regs$dump_out$007;
  assign snapshots$001$set_in_$008      = regs$dump_out$008;
  assign snapshots$001$set_in_$009      = regs$dump_out$009;
  assign snapshots$001$set_in_$010      = regs$dump_out$010;
  assign snapshots$001$set_in_$011      = regs$dump_out$011;
  assign snapshots$001$set_in_$012      = regs$dump_out$012;
  assign snapshots$001$set_in_$013      = regs$dump_out$013;
  assign snapshots$001$set_in_$014      = regs$dump_out$014;
  assign snapshots$001$set_in_$015      = regs$dump_out$015;
  assign snapshots$001$set_in_$016      = regs$dump_out$016;
  assign snapshots$001$set_in_$017      = regs$dump_out$017;
  assign snapshots$001$set_in_$018      = regs$dump_out$018;
  assign snapshots$001$set_in_$019      = regs$dump_out$019;
  assign snapshots$001$set_in_$020      = regs$dump_out$020;
  assign snapshots$001$set_in_$021      = regs$dump_out$021;
  assign snapshots$001$set_in_$022      = regs$dump_out$022;
  assign snapshots$001$set_in_$023      = regs$dump_out$023;
  assign snapshots$001$set_in_$024      = regs$dump_out$024;
  assign snapshots$001$set_in_$025      = regs$dump_out$025;
  assign snapshots$001$set_in_$026      = regs$dump_out$026;
  assign snapshots$001$set_in_$027      = regs$dump_out$027;
  assign snapshots$001$set_in_$028      = regs$dump_out$028;
  assign snapshots$001$set_in_$029      = regs$dump_out$029;
  assign snapshots$001$set_in_$030      = regs$dump_out$030;
  assign snapshots$001$set_in_$031      = regs$dump_out$031;

  // array declarations
  logic    [   0:0] snapshots$set_call[0:1];
  assign snapshots$000$set_call = snapshots$set_call[  0];
  assign snapshots$001$set_call = snapshots$set_call[  1];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_snapshot_save(i=i):
  //         s.snapshots[
  //             i].set_call.v = s.snapshot_call and s.snapshot_target_id == i

  // logic for handle_snapshot_save()
  always @ (*) begin
    snapshots$set_call[0] = (snapshot_call&&(snapshot_target_id == 0));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_snapshot_save(i=i):
  //         s.snapshots[
  //             i].set_call.v = s.snapshot_call and s.snapshot_target_id == i

  // logic for handle_snapshot_save()
  always @ (*) begin
    snapshots$set_call[1] = (snapshot_call&&(snapshot_target_id == 1));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_should_restore(j=j):
  //           if s.snapshot_call and s.restore_call and s.snapshot_target_id == s.restore_source_id:
  //             s.should_restore.v = 0
  //           else:
  //             s.should_restore.v = s.restore_call

  // logic for compute_should_restore()
  always @ (*) begin
    if ((snapshot_call&&restore_call&&(snapshot_target_id == restore_source_id))) begin
      should_restore = 0;
    end
    else begin
      should_restore = restore_call;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_should_set():
  //       s.should_set.v = s.should_restore | s.set_call

  // logic for handle_should_set()
  always @ (*) begin
    should_set = (should_restore|set_call);
  end


endmodule // SnapshottingRegisterFile_0x66bdadc3daaa062

//-----------------------------------------------------------------------------
// RegisterFile_0x7c767f76bd64c12c
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.registerfile {"dtype": 6, "nregs": 32, "num_read_ports": 2, "num_write_ports": 1, "reset_values": [0, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30], "write_dump_bypass": true, "write_read_bypass": false}
// PyMTL: verilator_xinit = zeros
module RegisterFile_0x7c767f76bd64c12c
(
  input  logic [   0:0] clk,
  output logic [   5:0] dump_out$000,
  output logic [   5:0] dump_out$010,
  output logic [   5:0] dump_out$011,
  output logic [   5:0] dump_out$012,
  output logic [   5:0] dump_out$013,
  output logic [   5:0] dump_out$014,
  output logic [   5:0] dump_out$015,
  output logic [   5:0] dump_out$016,
  output logic [   5:0] dump_out$017,
  output logic [   5:0] dump_out$018,
  output logic [   5:0] dump_out$019,
  output logic [   5:0] dump_out$001,
  output logic [   5:0] dump_out$020,
  output logic [   5:0] dump_out$021,
  output logic [   5:0] dump_out$022,
  output logic [   5:0] dump_out$023,
  output logic [   5:0] dump_out$024,
  output logic [   5:0] dump_out$025,
  output logic [   5:0] dump_out$026,
  output logic [   5:0] dump_out$027,
  output logic [   5:0] dump_out$028,
  output logic [   5:0] dump_out$029,
  output logic [   5:0] dump_out$002,
  output logic [   5:0] dump_out$030,
  output logic [   5:0] dump_out$031,
  output logic [   5:0] dump_out$003,
  output logic [   5:0] dump_out$004,
  output logic [   5:0] dump_out$005,
  output logic [   5:0] dump_out$006,
  output logic [   5:0] dump_out$007,
  output logic [   5:0] dump_out$008,
  output logic [   5:0] dump_out$009,
  input  logic [   4:0] read_addr$000,
  input  logic [   4:0] read_addr$001,
  output logic [   5:0] read_data$000,
  output logic [   5:0] read_data$001,
  input  logic [   0:0] reset,
  input  logic [   0:0] set_call,
  input  logic [   5:0] set_in_$000,
  input  logic [   5:0] set_in_$010,
  input  logic [   5:0] set_in_$011,
  input  logic [   5:0] set_in_$012,
  input  logic [   5:0] set_in_$013,
  input  logic [   5:0] set_in_$014,
  input  logic [   5:0] set_in_$015,
  input  logic [   5:0] set_in_$016,
  input  logic [   5:0] set_in_$017,
  input  logic [   5:0] set_in_$018,
  input  logic [   5:0] set_in_$019,
  input  logic [   5:0] set_in_$001,
  input  logic [   5:0] set_in_$020,
  input  logic [   5:0] set_in_$021,
  input  logic [   5:0] set_in_$022,
  input  logic [   5:0] set_in_$023,
  input  logic [   5:0] set_in_$024,
  input  logic [   5:0] set_in_$025,
  input  logic [   5:0] set_in_$026,
  input  logic [   5:0] set_in_$027,
  input  logic [   5:0] set_in_$028,
  input  logic [   5:0] set_in_$029,
  input  logic [   5:0] set_in_$002,
  input  logic [   5:0] set_in_$030,
  input  logic [   5:0] set_in_$031,
  input  logic [   5:0] set_in_$003,
  input  logic [   5:0] set_in_$004,
  input  logic [   5:0] set_in_$005,
  input  logic [   5:0] set_in_$006,
  input  logic [   5:0] set_in_$007,
  input  logic [   5:0] set_in_$008,
  input  logic [   5:0] set_in_$009,
  input  logic [   4:0] write_addr$000,
  input  logic [   0:0] write_call$000,
  input  logic [   5:0] write_data$000
);

  // logic declarations
  logic   [   5:0] write_inc$000;
  logic   [   5:0] write_inc$001;
  logic   [   5:0] write_inc$002;
  logic   [   5:0] write_inc$003;
  logic   [   5:0] write_inc$004;
  logic   [   5:0] write_inc$005;
  logic   [   5:0] write_inc$006;
  logic   [   5:0] write_inc$007;
  logic   [   5:0] write_inc$008;
  logic   [   5:0] write_inc$009;
  logic   [   5:0] write_inc$010;
  logic   [   5:0] write_inc$011;
  logic   [   5:0] write_inc$012;
  logic   [   5:0] write_inc$013;
  logic   [   5:0] write_inc$014;
  logic   [   5:0] write_inc$015;
  logic   [   5:0] write_inc$016;
  logic   [   5:0] write_inc$017;
  logic   [   5:0] write_inc$018;
  logic   [   5:0] write_inc$019;
  logic   [   5:0] write_inc$020;
  logic   [   5:0] write_inc$021;
  logic   [   5:0] write_inc$022;
  logic   [   5:0] write_inc$023;
  logic   [   5:0] write_inc$024;
  logic   [   5:0] write_inc$025;
  logic   [   5:0] write_inc$026;
  logic   [   5:0] write_inc$027;
  logic   [   5:0] write_inc$028;
  logic   [   5:0] write_inc$029;
  logic   [   5:0] write_inc$030;
  logic   [   5:0] write_inc$031;
  logic   [   5:0] after_set$000;
  logic   [   5:0] after_set$001;
  logic   [   5:0] after_set$002;
  logic   [   5:0] after_set$003;
  logic   [   5:0] after_set$004;
  logic   [   5:0] after_set$005;
  logic   [   5:0] after_set$006;
  logic   [   5:0] after_set$007;
  logic   [   5:0] after_set$008;
  logic   [   5:0] after_set$009;
  logic   [   5:0] after_set$010;
  logic   [   5:0] after_set$011;
  logic   [   5:0] after_set$012;
  logic   [   5:0] after_set$013;
  logic   [   5:0] after_set$014;
  logic   [   5:0] after_set$015;
  logic   [   5:0] after_set$016;
  logic   [   5:0] after_set$017;
  logic   [   5:0] after_set$018;
  logic   [   5:0] after_set$019;
  logic   [   5:0] after_set$020;
  logic   [   5:0] after_set$021;
  logic   [   5:0] after_set$022;
  logic   [   5:0] after_set$023;
  logic   [   5:0] after_set$024;
  logic   [   5:0] after_set$025;
  logic   [   5:0] after_set$026;
  logic   [   5:0] after_set$027;
  logic   [   5:0] after_set$028;
  logic   [   5:0] after_set$029;
  logic   [   5:0] after_set$030;
  logic   [   5:0] after_set$031;
  logic   [   5:0] regs$000;
  logic   [   5:0] regs$001;
  logic   [   5:0] regs$002;
  logic   [   5:0] regs$003;
  logic   [   5:0] regs$004;
  logic   [   5:0] regs$005;
  logic   [   5:0] regs$006;
  logic   [   5:0] regs$007;
  logic   [   5:0] regs$008;
  logic   [   5:0] regs$009;
  logic   [   5:0] regs$010;
  logic   [   5:0] regs$011;
  logic   [   5:0] regs$012;
  logic   [   5:0] regs$013;
  logic   [   5:0] regs$014;
  logic   [   5:0] regs$015;
  logic   [   5:0] regs$016;
  logic   [   5:0] regs$017;
  logic   [   5:0] regs$018;
  logic   [   5:0] regs$019;
  logic   [   5:0] regs$020;
  logic   [   5:0] regs$021;
  logic   [   5:0] regs$022;
  logic   [   5:0] regs$023;
  logic   [   5:0] regs$024;
  logic   [   5:0] regs$025;
  logic   [   5:0] regs$026;
  logic   [   5:0] regs$027;
  logic   [   5:0] regs$028;
  logic   [   5:0] regs$029;
  logic   [   5:0] regs$030;
  logic   [   5:0] regs$031;
  logic   [   5:0] after_write$000;
  logic   [   5:0] after_write$001;
  logic   [   5:0] after_write$002;
  logic   [   5:0] after_write$003;
  logic   [   5:0] after_write$004;
  logic   [   5:0] after_write$005;
  logic   [   5:0] after_write$006;
  logic   [   5:0] after_write$007;
  logic   [   5:0] after_write$008;
  logic   [   5:0] after_write$009;
  logic   [   5:0] after_write$010;
  logic   [   5:0] after_write$011;
  logic   [   5:0] after_write$012;
  logic   [   5:0] after_write$013;
  logic   [   5:0] after_write$014;
  logic   [   5:0] after_write$015;
  logic   [   5:0] after_write$016;
  logic   [   5:0] after_write$017;
  logic   [   5:0] after_write$018;
  logic   [   5:0] after_write$019;
  logic   [   5:0] after_write$020;
  logic   [   5:0] after_write$021;
  logic   [   5:0] after_write$022;
  logic   [   5:0] after_write$023;
  logic   [   5:0] after_write$024;
  logic   [   5:0] after_write$025;
  logic   [   5:0] after_write$026;
  logic   [   5:0] after_write$027;
  logic   [   5:0] after_write$028;
  logic   [   5:0] after_write$029;
  logic   [   5:0] after_write$030;
  logic   [   5:0] after_write$031;


  // signal connections
  assign dump_out$000 = after_write$000;
  assign dump_out$001 = after_write$001;
  assign dump_out$002 = after_write$002;
  assign dump_out$003 = after_write$003;
  assign dump_out$004 = after_write$004;
  assign dump_out$005 = after_write$005;
  assign dump_out$006 = after_write$006;
  assign dump_out$007 = after_write$007;
  assign dump_out$008 = after_write$008;
  assign dump_out$009 = after_write$009;
  assign dump_out$010 = after_write$010;
  assign dump_out$011 = after_write$011;
  assign dump_out$012 = after_write$012;
  assign dump_out$013 = after_write$013;
  assign dump_out$014 = after_write$014;
  assign dump_out$015 = after_write$015;
  assign dump_out$016 = after_write$016;
  assign dump_out$017 = after_write$017;
  assign dump_out$018 = after_write$018;
  assign dump_out$019 = after_write$019;
  assign dump_out$020 = after_write$020;
  assign dump_out$021 = after_write$021;
  assign dump_out$022 = after_write$022;
  assign dump_out$023 = after_write$023;
  assign dump_out$024 = after_write$024;
  assign dump_out$025 = after_write$025;
  assign dump_out$026 = after_write$026;
  assign dump_out$027 = after_write$027;
  assign dump_out$028 = after_write$028;
  assign dump_out$029 = after_write$029;
  assign dump_out$030 = after_write$030;
  assign dump_out$031 = after_write$031;

  // array declarations
  logic    [   5:0] after_set[0:31];
  assign after_set$000 = after_set[  0];
  assign after_set$001 = after_set[  1];
  assign after_set$002 = after_set[  2];
  assign after_set$003 = after_set[  3];
  assign after_set$004 = after_set[  4];
  assign after_set$005 = after_set[  5];
  assign after_set$006 = after_set[  6];
  assign after_set$007 = after_set[  7];
  assign after_set$008 = after_set[  8];
  assign after_set$009 = after_set[  9];
  assign after_set$010 = after_set[ 10];
  assign after_set$011 = after_set[ 11];
  assign after_set$012 = after_set[ 12];
  assign after_set$013 = after_set[ 13];
  assign after_set$014 = after_set[ 14];
  assign after_set$015 = after_set[ 15];
  assign after_set$016 = after_set[ 16];
  assign after_set$017 = after_set[ 17];
  assign after_set$018 = after_set[ 18];
  assign after_set$019 = after_set[ 19];
  assign after_set$020 = after_set[ 20];
  assign after_set$021 = after_set[ 21];
  assign after_set$022 = after_set[ 22];
  assign after_set$023 = after_set[ 23];
  assign after_set$024 = after_set[ 24];
  assign after_set$025 = after_set[ 25];
  assign after_set$026 = after_set[ 26];
  assign after_set$027 = after_set[ 27];
  assign after_set$028 = after_set[ 28];
  assign after_set$029 = after_set[ 29];
  assign after_set$030 = after_set[ 30];
  assign after_set$031 = after_set[ 31];
  logic    [   5:0] after_write[0:31];
  assign after_write$000 = after_write[  0];
  assign after_write$001 = after_write[  1];
  assign after_write$002 = after_write[  2];
  assign after_write$003 = after_write[  3];
  assign after_write$004 = after_write[  4];
  assign after_write$005 = after_write[  5];
  assign after_write$006 = after_write[  6];
  assign after_write$007 = after_write[  7];
  assign after_write$008 = after_write[  8];
  assign after_write$009 = after_write[  9];
  assign after_write$010 = after_write[ 10];
  assign after_write$011 = after_write[ 11];
  assign after_write$012 = after_write[ 12];
  assign after_write$013 = after_write[ 13];
  assign after_write$014 = after_write[ 14];
  assign after_write$015 = after_write[ 15];
  assign after_write$016 = after_write[ 16];
  assign after_write$017 = after_write[ 17];
  assign after_write$018 = after_write[ 18];
  assign after_write$019 = after_write[ 19];
  assign after_write$020 = after_write[ 20];
  assign after_write$021 = after_write[ 21];
  assign after_write$022 = after_write[ 22];
  assign after_write$023 = after_write[ 23];
  assign after_write$024 = after_write[ 24];
  assign after_write$025 = after_write[ 25];
  assign after_write$026 = after_write[ 26];
  assign after_write$027 = after_write[ 27];
  assign after_write$028 = after_write[ 28];
  assign after_write$029 = after_write[ 29];
  assign after_write$030 = after_write[ 30];
  assign after_write$031 = after_write[ 31];
  logic   [   4:0] read_addr[0:1];
  assign read_addr[  0] = read_addr$000;
  assign read_addr[  1] = read_addr$001;
  logic    [   5:0] read_data[0:1];
  assign read_data$000 = read_data[  0];
  assign read_data$001 = read_data[  1];
  logic    [   5:0] regs[0:31];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  assign regs$002 = regs[  2];
  assign regs$003 = regs[  3];
  assign regs$004 = regs[  4];
  assign regs$005 = regs[  5];
  assign regs$006 = regs[  6];
  assign regs$007 = regs[  7];
  assign regs$008 = regs[  8];
  assign regs$009 = regs[  9];
  assign regs$010 = regs[ 10];
  assign regs$011 = regs[ 11];
  assign regs$012 = regs[ 12];
  assign regs$013 = regs[ 13];
  assign regs$014 = regs[ 14];
  assign regs$015 = regs[ 15];
  assign regs$016 = regs[ 16];
  assign regs$017 = regs[ 17];
  assign regs$018 = regs[ 18];
  assign regs$019 = regs[ 19];
  assign regs$020 = regs[ 20];
  assign regs$021 = regs[ 21];
  assign regs$022 = regs[ 22];
  assign regs$023 = regs[ 23];
  assign regs$024 = regs[ 24];
  assign regs$025 = regs[ 25];
  assign regs$026 = regs[ 26];
  assign regs$027 = regs[ 27];
  assign regs$028 = regs[ 28];
  assign regs$029 = regs[ 29];
  assign regs$030 = regs[ 30];
  assign regs$031 = regs[ 31];
  logic   [   5:0] set_in_[0:31];
  assign set_in_[  0] = set_in_$000;
  assign set_in_[  1] = set_in_$001;
  assign set_in_[  2] = set_in_$002;
  assign set_in_[  3] = set_in_$003;
  assign set_in_[  4] = set_in_$004;
  assign set_in_[  5] = set_in_$005;
  assign set_in_[  6] = set_in_$006;
  assign set_in_[  7] = set_in_$007;
  assign set_in_[  8] = set_in_$008;
  assign set_in_[  9] = set_in_$009;
  assign set_in_[ 10] = set_in_$010;
  assign set_in_[ 11] = set_in_$011;
  assign set_in_[ 12] = set_in_$012;
  assign set_in_[ 13] = set_in_$013;
  assign set_in_[ 14] = set_in_$014;
  assign set_in_[ 15] = set_in_$015;
  assign set_in_[ 16] = set_in_$016;
  assign set_in_[ 17] = set_in_$017;
  assign set_in_[ 18] = set_in_$018;
  assign set_in_[ 19] = set_in_$019;
  assign set_in_[ 20] = set_in_$020;
  assign set_in_[ 21] = set_in_$021;
  assign set_in_[ 22] = set_in_$022;
  assign set_in_[ 23] = set_in_$023;
  assign set_in_[ 24] = set_in_$024;
  assign set_in_[ 25] = set_in_$025;
  assign set_in_[ 26] = set_in_$026;
  assign set_in_[ 27] = set_in_$027;
  assign set_in_[ 28] = set_in_$028;
  assign set_in_[ 29] = set_in_$029;
  assign set_in_[ 30] = set_in_$030;
  assign set_in_[ 31] = set_in_$031;
  logic   [   4:0] write_addr[0:0];
  assign write_addr[  0] = write_addr$000;
  logic   [   0:0] write_call[0:0];
  assign write_call[  0] = write_call$000;
  logic   [   5:0] write_data[0:0];
  assign write_data[  0] = write_data$000;
  logic    [   5:0] write_inc[0:31];
  assign write_inc$000 = write_inc[  0];
  assign write_inc$001 = write_inc[  1];
  assign write_inc$002 = write_inc[  2];
  assign write_inc$003 = write_inc[  3];
  assign write_inc$004 = write_inc[  4];
  assign write_inc$005 = write_inc[  5];
  assign write_inc$006 = write_inc[  6];
  assign write_inc$007 = write_inc[  7];
  assign write_inc$008 = write_inc[  8];
  assign write_inc$009 = write_inc[  9];
  assign write_inc$010 = write_inc[ 10];
  assign write_inc$011 = write_inc[ 11];
  assign write_inc$012 = write_inc[ 12];
  assign write_inc$013 = write_inc[ 13];
  assign write_inc$014 = write_inc[ 14];
  assign write_inc$015 = write_inc[ 15];
  assign write_inc$016 = write_inc[ 16];
  assign write_inc$017 = write_inc[ 17];
  assign write_inc$018 = write_inc[ 18];
  assign write_inc$019 = write_inc[ 19];
  assign write_inc$020 = write_inc[ 20];
  assign write_inc$021 = write_inc[ 21];
  assign write_inc$022 = write_inc[ 22];
  assign write_inc$023 = write_inc[ 23];
  assign write_inc$024 = write_inc[ 24];
  assign write_inc$025 = write_inc[ 25];
  assign write_inc$026 = write_inc[ 26];
  assign write_inc$027 = write_inc[ 27];
  assign write_inc$028 = write_inc[ 28];
  assign write_inc$029 = write_inc[ 29];
  assign write_inc$030 = write_inc[ 30];
  assign write_inc$031 = write_inc[ 31];

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[0] <= 0;
    end
    else begin
      regs[0] <= after_set[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[1] <= 0;
    end
    else begin
      regs[1] <= after_set[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[2] <= 1;
    end
    else begin
      regs[2] <= after_set[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[3] <= 2;
    end
    else begin
      regs[3] <= after_set[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[4] <= 3;
    end
    else begin
      regs[4] <= after_set[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[5] <= 4;
    end
    else begin
      regs[5] <= after_set[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[6] <= 5;
    end
    else begin
      regs[6] <= after_set[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[7] <= 6;
    end
    else begin
      regs[7] <= after_set[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[8] <= 7;
    end
    else begin
      regs[8] <= after_set[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[9] <= 8;
    end
    else begin
      regs[9] <= after_set[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[10] <= 9;
    end
    else begin
      regs[10] <= after_set[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[11] <= 10;
    end
    else begin
      regs[11] <= after_set[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[12] <= 11;
    end
    else begin
      regs[12] <= after_set[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[13] <= 12;
    end
    else begin
      regs[13] <= after_set[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[14] <= 13;
    end
    else begin
      regs[14] <= after_set[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[15] <= 14;
    end
    else begin
      regs[15] <= after_set[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[16] <= 15;
    end
    else begin
      regs[16] <= after_set[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[17] <= 16;
    end
    else begin
      regs[17] <= after_set[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[18] <= 17;
    end
    else begin
      regs[18] <= after_set[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[19] <= 18;
    end
    else begin
      regs[19] <= after_set[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[20] <= 19;
    end
    else begin
      regs[20] <= after_set[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[21] <= 20;
    end
    else begin
      regs[21] <= after_set[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[22] <= 21;
    end
    else begin
      regs[22] <= after_set[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[23] <= 22;
    end
    else begin
      regs[23] <= after_set[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[24] <= 23;
    end
    else begin
      regs[24] <= after_set[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[25] <= 24;
    end
    else begin
      regs[25] <= after_set[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[26] <= 25;
    end
    else begin
      regs[26] <= after_set[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[27] <= 26;
    end
    else begin
      regs[27] <= after_set[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[28] <= 27;
    end
    else begin
      regs[28] <= after_set[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[29] <= 28;
    end
    else begin
      regs[29] <= after_set[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[30] <= 29;
    end
    else begin
      regs[30] <= after_set[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[31] <= 30;
    end
    else begin
      regs[31] <= after_set[31];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 0))) begin
      write_inc[0] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[0] = regs[0];
      end
      else begin
        write_inc[0] = write_inc[-32];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[0] = write_inc[0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[0] = set_in_[0];
    end
    else begin
      after_set[0] = after_write[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 1))) begin
      write_inc[1] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[1] = regs[1];
      end
      else begin
        write_inc[1] = write_inc[-31];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[1] = write_inc[1];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[1] = set_in_[1];
    end
    else begin
      after_set[1] = after_write[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 2))) begin
      write_inc[2] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[2] = regs[2];
      end
      else begin
        write_inc[2] = write_inc[-30];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[2] = write_inc[2];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[2] = set_in_[2];
    end
    else begin
      after_set[2] = after_write[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 3))) begin
      write_inc[3] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[3] = regs[3];
      end
      else begin
        write_inc[3] = write_inc[-29];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[3] = write_inc[3];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[3] = set_in_[3];
    end
    else begin
      after_set[3] = after_write[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 4))) begin
      write_inc[4] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[4] = regs[4];
      end
      else begin
        write_inc[4] = write_inc[-28];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[4] = write_inc[4];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[4] = set_in_[4];
    end
    else begin
      after_set[4] = after_write[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 5))) begin
      write_inc[5] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[5] = regs[5];
      end
      else begin
        write_inc[5] = write_inc[-27];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[5] = write_inc[5];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[5] = set_in_[5];
    end
    else begin
      after_set[5] = after_write[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 6))) begin
      write_inc[6] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[6] = regs[6];
      end
      else begin
        write_inc[6] = write_inc[-26];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[6] = write_inc[6];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[6] = set_in_[6];
    end
    else begin
      after_set[6] = after_write[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 7))) begin
      write_inc[7] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[7] = regs[7];
      end
      else begin
        write_inc[7] = write_inc[-25];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[7] = write_inc[7];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[7] = set_in_[7];
    end
    else begin
      after_set[7] = after_write[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 8))) begin
      write_inc[8] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[8] = regs[8];
      end
      else begin
        write_inc[8] = write_inc[-24];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[8] = write_inc[8];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[8] = set_in_[8];
    end
    else begin
      after_set[8] = after_write[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 9))) begin
      write_inc[9] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[9] = regs[9];
      end
      else begin
        write_inc[9] = write_inc[-23];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[9] = write_inc[9];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[9] = set_in_[9];
    end
    else begin
      after_set[9] = after_write[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 10))) begin
      write_inc[10] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[10] = regs[10];
      end
      else begin
        write_inc[10] = write_inc[-22];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[10] = write_inc[10];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[10] = set_in_[10];
    end
    else begin
      after_set[10] = after_write[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 11))) begin
      write_inc[11] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[11] = regs[11];
      end
      else begin
        write_inc[11] = write_inc[-21];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[11] = write_inc[11];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[11] = set_in_[11];
    end
    else begin
      after_set[11] = after_write[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 12))) begin
      write_inc[12] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[12] = regs[12];
      end
      else begin
        write_inc[12] = write_inc[-20];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[12] = write_inc[12];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[12] = set_in_[12];
    end
    else begin
      after_set[12] = after_write[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 13))) begin
      write_inc[13] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[13] = regs[13];
      end
      else begin
        write_inc[13] = write_inc[-19];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[13] = write_inc[13];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[13] = set_in_[13];
    end
    else begin
      after_set[13] = after_write[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 14))) begin
      write_inc[14] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[14] = regs[14];
      end
      else begin
        write_inc[14] = write_inc[-18];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[14] = write_inc[14];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[14] = set_in_[14];
    end
    else begin
      after_set[14] = after_write[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 15))) begin
      write_inc[15] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[15] = regs[15];
      end
      else begin
        write_inc[15] = write_inc[-17];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[15] = write_inc[15];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[15] = set_in_[15];
    end
    else begin
      after_set[15] = after_write[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 16))) begin
      write_inc[16] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[16] = regs[16];
      end
      else begin
        write_inc[16] = write_inc[-16];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[16] = write_inc[16];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[16] = set_in_[16];
    end
    else begin
      after_set[16] = after_write[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 17))) begin
      write_inc[17] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[17] = regs[17];
      end
      else begin
        write_inc[17] = write_inc[-15];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[17] = write_inc[17];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[17] = set_in_[17];
    end
    else begin
      after_set[17] = after_write[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 18))) begin
      write_inc[18] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[18] = regs[18];
      end
      else begin
        write_inc[18] = write_inc[-14];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[18] = write_inc[18];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[18] = set_in_[18];
    end
    else begin
      after_set[18] = after_write[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 19))) begin
      write_inc[19] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[19] = regs[19];
      end
      else begin
        write_inc[19] = write_inc[-13];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[19] = write_inc[19];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[19] = set_in_[19];
    end
    else begin
      after_set[19] = after_write[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 20))) begin
      write_inc[20] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[20] = regs[20];
      end
      else begin
        write_inc[20] = write_inc[-12];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[20] = write_inc[20];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[20] = set_in_[20];
    end
    else begin
      after_set[20] = after_write[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 21))) begin
      write_inc[21] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[21] = regs[21];
      end
      else begin
        write_inc[21] = write_inc[-11];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[21] = write_inc[21];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[21] = set_in_[21];
    end
    else begin
      after_set[21] = after_write[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 22))) begin
      write_inc[22] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[22] = regs[22];
      end
      else begin
        write_inc[22] = write_inc[-10];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[22] = write_inc[22];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[22] = set_in_[22];
    end
    else begin
      after_set[22] = after_write[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 23))) begin
      write_inc[23] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[23] = regs[23];
      end
      else begin
        write_inc[23] = write_inc[-9];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[23] = write_inc[23];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[23] = set_in_[23];
    end
    else begin
      after_set[23] = after_write[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 24))) begin
      write_inc[24] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[24] = regs[24];
      end
      else begin
        write_inc[24] = write_inc[-8];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[24] = write_inc[24];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[24] = set_in_[24];
    end
    else begin
      after_set[24] = after_write[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 25))) begin
      write_inc[25] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[25] = regs[25];
      end
      else begin
        write_inc[25] = write_inc[-7];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[25] = write_inc[25];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[25] = set_in_[25];
    end
    else begin
      after_set[25] = after_write[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 26))) begin
      write_inc[26] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[26] = regs[26];
      end
      else begin
        write_inc[26] = write_inc[-6];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[26] = write_inc[26];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[26] = set_in_[26];
    end
    else begin
      after_set[26] = after_write[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 27))) begin
      write_inc[27] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[27] = regs[27];
      end
      else begin
        write_inc[27] = write_inc[-5];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[27] = write_inc[27];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[27] = set_in_[27];
    end
    else begin
      after_set[27] = after_write[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 28))) begin
      write_inc[28] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[28] = regs[28];
      end
      else begin
        write_inc[28] = write_inc[-4];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[28] = write_inc[28];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[28] = set_in_[28];
    end
    else begin
      after_set[28] = after_write[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 29))) begin
      write_inc[29] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[29] = regs[29];
      end
      else begin
        write_inc[29] = write_inc[-3];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[29] = write_inc[29];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[29] = set_in_[29];
    end
    else begin
      after_set[29] = after_write[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 30))) begin
      write_inc[30] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[30] = regs[30];
      end
      else begin
        write_inc[30] = write_inc[-2];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[30] = write_inc[30];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[30] = set_in_[30];
    end
    else begin
      after_set[30] = after_write[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 31))) begin
      write_inc[31] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[31] = regs[31];
      end
      else begin
        write_inc[31] = write_inc[-1];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[31] = write_inc[31];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[31] = set_in_[31];
    end
    else begin
      after_set[31] = after_write[31];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_read(port=port):
  //           s.read_data[port].v = s.regs[s.read_addr[port]]

  // logic for handle_read()
  always @ (*) begin
    read_data[0] = regs[read_addr[0]];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_read(port=port):
  //           s.read_data[port].v = s.regs[s.read_addr[port]]

  // logic for handle_read()
  always @ (*) begin
    read_data[1] = regs[read_addr[1]];
  end


endmodule // RegisterFile_0x7c767f76bd64c12c

//-----------------------------------------------------------------------------
// Mux_0x387678144da2c8e
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.mux {"dtype": 6, "nports": 2}
// PyMTL: verilator_xinit = zeros
module Mux_0x387678144da2c8e
(
  input  logic [   0:0] clk,
  input  logic [   5:0] mux_in_$000,
  input  logic [   5:0] mux_in_$001,
  output logic  [   5:0] mux_out,
  input  logic [   0:0] mux_select,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nports = 2;


  // array declarations
  logic   [   5:0] mux_in_[0:1];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def select():
  //       assert s.mux_select < nports
  //       s.mux_out.v = s.mux_in_[s.mux_select]

  // logic for select()
  always @ (*) begin
    mux_out = mux_in_[mux_select];
  end


endmodule // Mux_0x387678144da2c8e

//-----------------------------------------------------------------------------
// RegisterFile_0x5b973c72ce6092d
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.registerfile {"dtype": 6, "nregs": 32, "num_read_ports": 0, "num_write_ports": 0, "reset_values": null, "write_dump_bypass": false, "write_read_bypass": false}
// PyMTL: verilator_xinit = zeros
module RegisterFile_0x5b973c72ce6092d
(
  input  logic [   0:0] clk,
  output logic [   5:0] dump_out$000,
  output logic [   5:0] dump_out$010,
  output logic [   5:0] dump_out$011,
  output logic [   5:0] dump_out$012,
  output logic [   5:0] dump_out$013,
  output logic [   5:0] dump_out$014,
  output logic [   5:0] dump_out$015,
  output logic [   5:0] dump_out$016,
  output logic [   5:0] dump_out$017,
  output logic [   5:0] dump_out$018,
  output logic [   5:0] dump_out$019,
  output logic [   5:0] dump_out$001,
  output logic [   5:0] dump_out$020,
  output logic [   5:0] dump_out$021,
  output logic [   5:0] dump_out$022,
  output logic [   5:0] dump_out$023,
  output logic [   5:0] dump_out$024,
  output logic [   5:0] dump_out$025,
  output logic [   5:0] dump_out$026,
  output logic [   5:0] dump_out$027,
  output logic [   5:0] dump_out$028,
  output logic [   5:0] dump_out$029,
  output logic [   5:0] dump_out$002,
  output logic [   5:0] dump_out$030,
  output logic [   5:0] dump_out$031,
  output logic [   5:0] dump_out$003,
  output logic [   5:0] dump_out$004,
  output logic [   5:0] dump_out$005,
  output logic [   5:0] dump_out$006,
  output logic [   5:0] dump_out$007,
  output logic [   5:0] dump_out$008,
  output logic [   5:0] dump_out$009,
  input  logic [   0:0] reset,
  input  logic [   0:0] set_call,
  input  logic [   5:0] set_in_$000,
  input  logic [   5:0] set_in_$010,
  input  logic [   5:0] set_in_$011,
  input  logic [   5:0] set_in_$012,
  input  logic [   5:0] set_in_$013,
  input  logic [   5:0] set_in_$014,
  input  logic [   5:0] set_in_$015,
  input  logic [   5:0] set_in_$016,
  input  logic [   5:0] set_in_$017,
  input  logic [   5:0] set_in_$018,
  input  logic [   5:0] set_in_$019,
  input  logic [   5:0] set_in_$001,
  input  logic [   5:0] set_in_$020,
  input  logic [   5:0] set_in_$021,
  input  logic [   5:0] set_in_$022,
  input  logic [   5:0] set_in_$023,
  input  logic [   5:0] set_in_$024,
  input  logic [   5:0] set_in_$025,
  input  logic [   5:0] set_in_$026,
  input  logic [   5:0] set_in_$027,
  input  logic [   5:0] set_in_$028,
  input  logic [   5:0] set_in_$029,
  input  logic [   5:0] set_in_$002,
  input  logic [   5:0] set_in_$030,
  input  logic [   5:0] set_in_$031,
  input  logic [   5:0] set_in_$003,
  input  logic [   5:0] set_in_$004,
  input  logic [   5:0] set_in_$005,
  input  logic [   5:0] set_in_$006,
  input  logic [   5:0] set_in_$007,
  input  logic [   5:0] set_in_$008,
  input  logic [   5:0] set_in_$009
);

  // logic declarations
  logic   [   5:0] after_set$000;
  logic   [   5:0] after_set$001;
  logic   [   5:0] after_set$002;
  logic   [   5:0] after_set$003;
  logic   [   5:0] after_set$004;
  logic   [   5:0] after_set$005;
  logic   [   5:0] after_set$006;
  logic   [   5:0] after_set$007;
  logic   [   5:0] after_set$008;
  logic   [   5:0] after_set$009;
  logic   [   5:0] after_set$010;
  logic   [   5:0] after_set$011;
  logic   [   5:0] after_set$012;
  logic   [   5:0] after_set$013;
  logic   [   5:0] after_set$014;
  logic   [   5:0] after_set$015;
  logic   [   5:0] after_set$016;
  logic   [   5:0] after_set$017;
  logic   [   5:0] after_set$018;
  logic   [   5:0] after_set$019;
  logic   [   5:0] after_set$020;
  logic   [   5:0] after_set$021;
  logic   [   5:0] after_set$022;
  logic   [   5:0] after_set$023;
  logic   [   5:0] after_set$024;
  logic   [   5:0] after_set$025;
  logic   [   5:0] after_set$026;
  logic   [   5:0] after_set$027;
  logic   [   5:0] after_set$028;
  logic   [   5:0] after_set$029;
  logic   [   5:0] after_set$030;
  logic   [   5:0] after_set$031;
  logic   [   5:0] regs$000;
  logic   [   5:0] regs$001;
  logic   [   5:0] regs$002;
  logic   [   5:0] regs$003;
  logic   [   5:0] regs$004;
  logic   [   5:0] regs$005;
  logic   [   5:0] regs$006;
  logic   [   5:0] regs$007;
  logic   [   5:0] regs$008;
  logic   [   5:0] regs$009;
  logic   [   5:0] regs$010;
  logic   [   5:0] regs$011;
  logic   [   5:0] regs$012;
  logic   [   5:0] regs$013;
  logic   [   5:0] regs$014;
  logic   [   5:0] regs$015;
  logic   [   5:0] regs$016;
  logic   [   5:0] regs$017;
  logic   [   5:0] regs$018;
  logic   [   5:0] regs$019;
  logic   [   5:0] regs$020;
  logic   [   5:0] regs$021;
  logic   [   5:0] regs$022;
  logic   [   5:0] regs$023;
  logic   [   5:0] regs$024;
  logic   [   5:0] regs$025;
  logic   [   5:0] regs$026;
  logic   [   5:0] regs$027;
  logic   [   5:0] regs$028;
  logic   [   5:0] regs$029;
  logic   [   5:0] regs$030;
  logic   [   5:0] regs$031;
  logic   [   5:0] after_write$000;
  logic   [   5:0] after_write$001;
  logic   [   5:0] after_write$002;
  logic   [   5:0] after_write$003;
  logic   [   5:0] after_write$004;
  logic   [   5:0] after_write$005;
  logic   [   5:0] after_write$006;
  logic   [   5:0] after_write$007;
  logic   [   5:0] after_write$008;
  logic   [   5:0] after_write$009;
  logic   [   5:0] after_write$010;
  logic   [   5:0] after_write$011;
  logic   [   5:0] after_write$012;
  logic   [   5:0] after_write$013;
  logic   [   5:0] after_write$014;
  logic   [   5:0] after_write$015;
  logic   [   5:0] after_write$016;
  logic   [   5:0] after_write$017;
  logic   [   5:0] after_write$018;
  logic   [   5:0] after_write$019;
  logic   [   5:0] after_write$020;
  logic   [   5:0] after_write$021;
  logic   [   5:0] after_write$022;
  logic   [   5:0] after_write$023;
  logic   [   5:0] after_write$024;
  logic   [   5:0] after_write$025;
  logic   [   5:0] after_write$026;
  logic   [   5:0] after_write$027;
  logic   [   5:0] after_write$028;
  logic   [   5:0] after_write$029;
  logic   [   5:0] after_write$030;
  logic   [   5:0] after_write$031;


  // signal connections
  assign dump_out$000 = regs$000;
  assign dump_out$001 = regs$001;
  assign dump_out$002 = regs$002;
  assign dump_out$003 = regs$003;
  assign dump_out$004 = regs$004;
  assign dump_out$005 = regs$005;
  assign dump_out$006 = regs$006;
  assign dump_out$007 = regs$007;
  assign dump_out$008 = regs$008;
  assign dump_out$009 = regs$009;
  assign dump_out$010 = regs$010;
  assign dump_out$011 = regs$011;
  assign dump_out$012 = regs$012;
  assign dump_out$013 = regs$013;
  assign dump_out$014 = regs$014;
  assign dump_out$015 = regs$015;
  assign dump_out$016 = regs$016;
  assign dump_out$017 = regs$017;
  assign dump_out$018 = regs$018;
  assign dump_out$019 = regs$019;
  assign dump_out$020 = regs$020;
  assign dump_out$021 = regs$021;
  assign dump_out$022 = regs$022;
  assign dump_out$023 = regs$023;
  assign dump_out$024 = regs$024;
  assign dump_out$025 = regs$025;
  assign dump_out$026 = regs$026;
  assign dump_out$027 = regs$027;
  assign dump_out$028 = regs$028;
  assign dump_out$029 = regs$029;
  assign dump_out$030 = regs$030;
  assign dump_out$031 = regs$031;

  // array declarations
  logic    [   5:0] after_set[0:31];
  assign after_set$000 = after_set[  0];
  assign after_set$001 = after_set[  1];
  assign after_set$002 = after_set[  2];
  assign after_set$003 = after_set[  3];
  assign after_set$004 = after_set[  4];
  assign after_set$005 = after_set[  5];
  assign after_set$006 = after_set[  6];
  assign after_set$007 = after_set[  7];
  assign after_set$008 = after_set[  8];
  assign after_set$009 = after_set[  9];
  assign after_set$010 = after_set[ 10];
  assign after_set$011 = after_set[ 11];
  assign after_set$012 = after_set[ 12];
  assign after_set$013 = after_set[ 13];
  assign after_set$014 = after_set[ 14];
  assign after_set$015 = after_set[ 15];
  assign after_set$016 = after_set[ 16];
  assign after_set$017 = after_set[ 17];
  assign after_set$018 = after_set[ 18];
  assign after_set$019 = after_set[ 19];
  assign after_set$020 = after_set[ 20];
  assign after_set$021 = after_set[ 21];
  assign after_set$022 = after_set[ 22];
  assign after_set$023 = after_set[ 23];
  assign after_set$024 = after_set[ 24];
  assign after_set$025 = after_set[ 25];
  assign after_set$026 = after_set[ 26];
  assign after_set$027 = after_set[ 27];
  assign after_set$028 = after_set[ 28];
  assign after_set$029 = after_set[ 29];
  assign after_set$030 = after_set[ 30];
  assign after_set$031 = after_set[ 31];
  logic    [   5:0] after_write[0:31];
  assign after_write$000 = after_write[  0];
  assign after_write$001 = after_write[  1];
  assign after_write$002 = after_write[  2];
  assign after_write$003 = after_write[  3];
  assign after_write$004 = after_write[  4];
  assign after_write$005 = after_write[  5];
  assign after_write$006 = after_write[  6];
  assign after_write$007 = after_write[  7];
  assign after_write$008 = after_write[  8];
  assign after_write$009 = after_write[  9];
  assign after_write$010 = after_write[ 10];
  assign after_write$011 = after_write[ 11];
  assign after_write$012 = after_write[ 12];
  assign after_write$013 = after_write[ 13];
  assign after_write$014 = after_write[ 14];
  assign after_write$015 = after_write[ 15];
  assign after_write$016 = after_write[ 16];
  assign after_write$017 = after_write[ 17];
  assign after_write$018 = after_write[ 18];
  assign after_write$019 = after_write[ 19];
  assign after_write$020 = after_write[ 20];
  assign after_write$021 = after_write[ 21];
  assign after_write$022 = after_write[ 22];
  assign after_write$023 = after_write[ 23];
  assign after_write$024 = after_write[ 24];
  assign after_write$025 = after_write[ 25];
  assign after_write$026 = after_write[ 26];
  assign after_write$027 = after_write[ 27];
  assign after_write$028 = after_write[ 28];
  assign after_write$029 = after_write[ 29];
  assign after_write$030 = after_write[ 30];
  assign after_write$031 = after_write[ 31];
  logic    [   5:0] regs[0:31];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  assign regs$002 = regs[  2];
  assign regs$003 = regs[  3];
  assign regs$004 = regs[  4];
  assign regs$005 = regs[  5];
  assign regs$006 = regs[  6];
  assign regs$007 = regs[  7];
  assign regs$008 = regs[  8];
  assign regs$009 = regs[  9];
  assign regs$010 = regs[ 10];
  assign regs$011 = regs[ 11];
  assign regs$012 = regs[ 12];
  assign regs$013 = regs[ 13];
  assign regs$014 = regs[ 14];
  assign regs$015 = regs[ 15];
  assign regs$016 = regs[ 16];
  assign regs$017 = regs[ 17];
  assign regs$018 = regs[ 18];
  assign regs$019 = regs[ 19];
  assign regs$020 = regs[ 20];
  assign regs$021 = regs[ 21];
  assign regs$022 = regs[ 22];
  assign regs$023 = regs[ 23];
  assign regs$024 = regs[ 24];
  assign regs$025 = regs[ 25];
  assign regs$026 = regs[ 26];
  assign regs$027 = regs[ 27];
  assign regs$028 = regs[ 28];
  assign regs$029 = regs[ 29];
  assign regs$030 = regs[ 30];
  assign regs$031 = regs[ 31];
  logic   [   5:0] set_in_[0:31];
  assign set_in_[  0] = set_in_$000;
  assign set_in_[  1] = set_in_$001;
  assign set_in_[  2] = set_in_$002;
  assign set_in_[  3] = set_in_$003;
  assign set_in_[  4] = set_in_$004;
  assign set_in_[  5] = set_in_$005;
  assign set_in_[  6] = set_in_$006;
  assign set_in_[  7] = set_in_$007;
  assign set_in_[  8] = set_in_$008;
  assign set_in_[  9] = set_in_$009;
  assign set_in_[ 10] = set_in_$010;
  assign set_in_[ 11] = set_in_$011;
  assign set_in_[ 12] = set_in_$012;
  assign set_in_[ 13] = set_in_$013;
  assign set_in_[ 14] = set_in_$014;
  assign set_in_[ 15] = set_in_$015;
  assign set_in_[ 16] = set_in_$016;
  assign set_in_[ 17] = set_in_$017;
  assign set_in_[ 18] = set_in_$018;
  assign set_in_[ 19] = set_in_$019;
  assign set_in_[ 20] = set_in_$020;
  assign set_in_[ 21] = set_in_$021;
  assign set_in_[ 22] = set_in_$022;
  assign set_in_[ 23] = set_in_$023;
  assign set_in_[ 24] = set_in_$024;
  assign set_in_[ 25] = set_in_$025;
  assign set_in_[ 26] = set_in_$026;
  assign set_in_[ 27] = set_in_$027;
  assign set_in_[ 28] = set_in_$028;
  assign set_in_[ 29] = set_in_$029;
  assign set_in_[ 30] = set_in_$030;
  assign set_in_[ 31] = set_in_$031;

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[0] <= 0;
    end
    else begin
      regs[0] <= after_set[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[1] <= 0;
    end
    else begin
      regs[1] <= after_set[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[2] <= 0;
    end
    else begin
      regs[2] <= after_set[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[3] <= 0;
    end
    else begin
      regs[3] <= after_set[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[4] <= 0;
    end
    else begin
      regs[4] <= after_set[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[5] <= 0;
    end
    else begin
      regs[5] <= after_set[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[6] <= 0;
    end
    else begin
      regs[6] <= after_set[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[7] <= 0;
    end
    else begin
      regs[7] <= after_set[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[8] <= 0;
    end
    else begin
      regs[8] <= after_set[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[9] <= 0;
    end
    else begin
      regs[9] <= after_set[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[10] <= 0;
    end
    else begin
      regs[10] <= after_set[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[11] <= 0;
    end
    else begin
      regs[11] <= after_set[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[12] <= 0;
    end
    else begin
      regs[12] <= after_set[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[13] <= 0;
    end
    else begin
      regs[13] <= after_set[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[14] <= 0;
    end
    else begin
      regs[14] <= after_set[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[15] <= 0;
    end
    else begin
      regs[15] <= after_set[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[16] <= 0;
    end
    else begin
      regs[16] <= after_set[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[17] <= 0;
    end
    else begin
      regs[17] <= after_set[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[18] <= 0;
    end
    else begin
      regs[18] <= after_set[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[19] <= 0;
    end
    else begin
      regs[19] <= after_set[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[20] <= 0;
    end
    else begin
      regs[20] <= after_set[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[21] <= 0;
    end
    else begin
      regs[21] <= after_set[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[22] <= 0;
    end
    else begin
      regs[22] <= after_set[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[23] <= 0;
    end
    else begin
      regs[23] <= after_set[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[24] <= 0;
    end
    else begin
      regs[24] <= after_set[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[25] <= 0;
    end
    else begin
      regs[25] <= after_set[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[26] <= 0;
    end
    else begin
      regs[26] <= after_set[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[27] <= 0;
    end
    else begin
      regs[27] <= after_set[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[28] <= 0;
    end
    else begin
      regs[28] <= after_set[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[29] <= 0;
    end
    else begin
      regs[29] <= after_set[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[30] <= 0;
    end
    else begin
      regs[30] <= after_set[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[31] <= 0;
    end
    else begin
      regs[31] <= after_set[31];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[0] = regs[0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[0] = set_in_[0];
    end
    else begin
      after_set[0] = after_write[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[1] = regs[1];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[1] = set_in_[1];
    end
    else begin
      after_set[1] = after_write[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[2] = regs[2];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[2] = set_in_[2];
    end
    else begin
      after_set[2] = after_write[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[3] = regs[3];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[3] = set_in_[3];
    end
    else begin
      after_set[3] = after_write[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[4] = regs[4];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[4] = set_in_[4];
    end
    else begin
      after_set[4] = after_write[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[5] = regs[5];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[5] = set_in_[5];
    end
    else begin
      after_set[5] = after_write[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[6] = regs[6];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[6] = set_in_[6];
    end
    else begin
      after_set[6] = after_write[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[7] = regs[7];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[7] = set_in_[7];
    end
    else begin
      after_set[7] = after_write[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[8] = regs[8];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[8] = set_in_[8];
    end
    else begin
      after_set[8] = after_write[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[9] = regs[9];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[9] = set_in_[9];
    end
    else begin
      after_set[9] = after_write[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[10] = regs[10];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[10] = set_in_[10];
    end
    else begin
      after_set[10] = after_write[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[11] = regs[11];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[11] = set_in_[11];
    end
    else begin
      after_set[11] = after_write[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[12] = regs[12];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[12] = set_in_[12];
    end
    else begin
      after_set[12] = after_write[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[13] = regs[13];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[13] = set_in_[13];
    end
    else begin
      after_set[13] = after_write[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[14] = regs[14];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[14] = set_in_[14];
    end
    else begin
      after_set[14] = after_write[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[15] = regs[15];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[15] = set_in_[15];
    end
    else begin
      after_set[15] = after_write[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[16] = regs[16];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[16] = set_in_[16];
    end
    else begin
      after_set[16] = after_write[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[17] = regs[17];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[17] = set_in_[17];
    end
    else begin
      after_set[17] = after_write[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[18] = regs[18];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[18] = set_in_[18];
    end
    else begin
      after_set[18] = after_write[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[19] = regs[19];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[19] = set_in_[19];
    end
    else begin
      after_set[19] = after_write[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[20] = regs[20];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[20] = set_in_[20];
    end
    else begin
      after_set[20] = after_write[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[21] = regs[21];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[21] = set_in_[21];
    end
    else begin
      after_set[21] = after_write[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[22] = regs[22];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[22] = set_in_[22];
    end
    else begin
      after_set[22] = after_write[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[23] = regs[23];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[23] = set_in_[23];
    end
    else begin
      after_set[23] = after_write[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[24] = regs[24];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[24] = set_in_[24];
    end
    else begin
      after_set[24] = after_write[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[25] = regs[25];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[25] = set_in_[25];
    end
    else begin
      after_set[25] = after_write[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[26] = regs[26];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[26] = set_in_[26];
    end
    else begin
      after_set[26] = after_write[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[27] = regs[27];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[27] = set_in_[27];
    end
    else begin
      after_set[27] = after_write[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[28] = regs[28];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[28] = set_in_[28];
    end
    else begin
      after_set[28] = after_write[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[29] = regs[29];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[29] = set_in_[29];
    end
    else begin
      after_set[29] = after_write[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[30] = regs[30];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[30] = set_in_[30];
    end
    else begin
      after_set[30] = after_write[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i):
  //           s.after_write[reg_i].v = s.regs[reg_i]

  // logic for update_last()
  always @ (*) begin
    after_write[31] = regs[31];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[31] = set_in_[31];
    end
    else begin
      after_set[31] = after_write[31];
    end
  end


endmodule // RegisterFile_0x5b973c72ce6092d

//-----------------------------------------------------------------------------
// AsynchronousRAM_0x6ff7d20a35694d13
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.async_ram {"interface": "write[1] <C> (data: Bits(5), addr: Bits(6)) -> (); read[1] (addr: Bits(6)) -> (data: Bits(5))", "reset_values": [1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00"]}
// PyMTL: verilator_xinit = zeros
module AsynchronousRAM_0x6ff7d20a35694d13
(
  input  logic [   0:0] clk,
  input  logic [   5:0] read_addr$000,
  output logic [   4:0] read_data$000,
  input  logic [   0:0] reset,
  input  logic [   5:0] write_addr$000,
  input  logic [   0:0] write_call$000,
  input  logic [   4:0] write_data$000
);

  // logic declarations
  logic   [   4:0] reset_values$000;
  logic   [   4:0] reset_values$001;
  logic   [   4:0] reset_values$002;
  logic   [   4:0] reset_values$003;
  logic   [   4:0] reset_values$004;
  logic   [   4:0] reset_values$005;
  logic   [   4:0] reset_values$006;
  logic   [   4:0] reset_values$007;
  logic   [   4:0] reset_values$008;
  logic   [   4:0] reset_values$009;
  logic   [   4:0] reset_values$010;
  logic   [   4:0] reset_values$011;
  logic   [   4:0] reset_values$012;
  logic   [   4:0] reset_values$013;
  logic   [   4:0] reset_values$014;
  logic   [   4:0] reset_values$015;
  logic   [   4:0] reset_values$016;
  logic   [   4:0] reset_values$017;
  logic   [   4:0] reset_values$018;
  logic   [   4:0] reset_values$019;
  logic   [   4:0] reset_values$020;
  logic   [   4:0] reset_values$021;
  logic   [   4:0] reset_values$022;
  logic   [   4:0] reset_values$023;
  logic   [   4:0] reset_values$024;
  logic   [   4:0] reset_values$025;
  logic   [   4:0] reset_values$026;
  logic   [   4:0] reset_values$027;
  logic   [   4:0] reset_values$028;
  logic   [   4:0] reset_values$029;
  logic   [   4:0] reset_values$030;
  logic   [   4:0] reset_values$031;
  logic   [   4:0] reset_values$032;
  logic   [   4:0] reset_values$033;
  logic   [   4:0] reset_values$034;
  logic   [   4:0] reset_values$035;
  logic   [   4:0] reset_values$036;
  logic   [   4:0] reset_values$037;
  logic   [   4:0] reset_values$038;
  logic   [   4:0] reset_values$039;
  logic   [   4:0] reset_values$040;
  logic   [   4:0] reset_values$041;
  logic   [   4:0] reset_values$042;
  logic   [   4:0] reset_values$043;
  logic   [   4:0] reset_values$044;
  logic   [   4:0] reset_values$045;
  logic   [   4:0] reset_values$046;
  logic   [   4:0] reset_values$047;
  logic   [   4:0] reset_values$048;
  logic   [   4:0] reset_values$049;
  logic   [   4:0] reset_values$050;
  logic   [   4:0] reset_values$051;
  logic   [   4:0] reset_values$052;
  logic   [   4:0] reset_values$053;
  logic   [   4:0] reset_values$054;
  logic   [   4:0] reset_values$055;
  logic   [   4:0] reset_values$056;
  logic   [   4:0] reset_values$057;
  logic   [   4:0] reset_values$058;
  logic   [   4:0] reset_values$059;
  logic   [   4:0] reset_values$060;
  logic   [   4:0] reset_values$061;
  logic   [   4:0] reset_values$062;
  logic   [   4:0] reset_values$063;
  logic   [   4:0] regs$000;
  logic   [   4:0] regs$001;
  logic   [   4:0] regs$002;
  logic   [   4:0] regs$003;
  logic   [   4:0] regs$004;
  logic   [   4:0] regs$005;
  logic   [   4:0] regs$006;
  logic   [   4:0] regs$007;
  logic   [   4:0] regs$008;
  logic   [   4:0] regs$009;
  logic   [   4:0] regs$010;
  logic   [   4:0] regs$011;
  logic   [   4:0] regs$012;
  logic   [   4:0] regs$013;
  logic   [   4:0] regs$014;
  logic   [   4:0] regs$015;
  logic   [   4:0] regs$016;
  logic   [   4:0] regs$017;
  logic   [   4:0] regs$018;
  logic   [   4:0] regs$019;
  logic   [   4:0] regs$020;
  logic   [   4:0] regs$021;
  logic   [   4:0] regs$022;
  logic   [   4:0] regs$023;
  logic   [   4:0] regs$024;
  logic   [   4:0] regs$025;
  logic   [   4:0] regs$026;
  logic   [   4:0] regs$027;
  logic   [   4:0] regs$028;
  logic   [   4:0] regs$029;
  logic   [   4:0] regs$030;
  logic   [   4:0] regs$031;
  logic   [   4:0] regs$032;
  logic   [   4:0] regs$033;
  logic   [   4:0] regs$034;
  logic   [   4:0] regs$035;
  logic   [   4:0] regs$036;
  logic   [   4:0] regs$037;
  logic   [   4:0] regs$038;
  logic   [   4:0] regs$039;
  logic   [   4:0] regs$040;
  logic   [   4:0] regs$041;
  logic   [   4:0] regs$042;
  logic   [   4:0] regs$043;
  logic   [   4:0] regs$044;
  logic   [   4:0] regs$045;
  logic   [   4:0] regs$046;
  logic   [   4:0] regs$047;
  logic   [   4:0] regs$048;
  logic   [   4:0] regs$049;
  logic   [   4:0] regs$050;
  logic   [   4:0] regs$051;
  logic   [   4:0] regs$052;
  logic   [   4:0] regs$053;
  logic   [   4:0] regs$054;
  logic   [   4:0] regs$055;
  logic   [   4:0] regs$056;
  logic   [   4:0] regs$057;
  logic   [   4:0] regs$058;
  logic   [   4:0] regs$059;
  logic   [   4:0] regs$060;
  logic   [   4:0] regs$061;
  logic   [   4:0] regs$062;
  logic   [   4:0] regs$063;


  // localparam declarations
  localparam num_read_ports = 1;
  localparam num_write_ports = 1;
  localparam nwords = 64;

  // loop variable declarations
  integer i;
  integer j;

  // signal connections
  assign reset_values$000 = 5'd1;
  assign reset_values$001 = 5'd2;
  assign reset_values$002 = 5'd3;
  assign reset_values$003 = 5'd4;
  assign reset_values$004 = 5'd5;
  assign reset_values$005 = 5'd6;
  assign reset_values$006 = 5'd7;
  assign reset_values$007 = 5'd8;
  assign reset_values$008 = 5'd9;
  assign reset_values$009 = 5'd10;
  assign reset_values$010 = 5'd11;
  assign reset_values$011 = 5'd12;
  assign reset_values$012 = 5'd13;
  assign reset_values$013 = 5'd14;
  assign reset_values$014 = 5'd15;
  assign reset_values$015 = 5'd16;
  assign reset_values$016 = 5'd17;
  assign reset_values$017 = 5'd18;
  assign reset_values$018 = 5'd19;
  assign reset_values$019 = 5'd20;
  assign reset_values$020 = 5'd21;
  assign reset_values$021 = 5'd22;
  assign reset_values$022 = 5'd23;
  assign reset_values$023 = 5'd24;
  assign reset_values$024 = 5'd25;
  assign reset_values$025 = 5'd26;
  assign reset_values$026 = 5'd27;
  assign reset_values$027 = 5'd28;
  assign reset_values$028 = 5'd29;
  assign reset_values$029 = 5'd30;
  assign reset_values$030 = 5'd31;
  assign reset_values$031 = 5'd0;
  assign reset_values$032 = 5'd0;
  assign reset_values$033 = 5'd0;
  assign reset_values$034 = 5'd0;
  assign reset_values$035 = 5'd0;
  assign reset_values$036 = 5'd0;
  assign reset_values$037 = 5'd0;
  assign reset_values$038 = 5'd0;
  assign reset_values$039 = 5'd0;
  assign reset_values$040 = 5'd0;
  assign reset_values$041 = 5'd0;
  assign reset_values$042 = 5'd0;
  assign reset_values$043 = 5'd0;
  assign reset_values$044 = 5'd0;
  assign reset_values$045 = 5'd0;
  assign reset_values$046 = 5'd0;
  assign reset_values$047 = 5'd0;
  assign reset_values$048 = 5'd0;
  assign reset_values$049 = 5'd0;
  assign reset_values$050 = 5'd0;
  assign reset_values$051 = 5'd0;
  assign reset_values$052 = 5'd0;
  assign reset_values$053 = 5'd0;
  assign reset_values$054 = 5'd0;
  assign reset_values$055 = 5'd0;
  assign reset_values$056 = 5'd0;
  assign reset_values$057 = 5'd0;
  assign reset_values$058 = 5'd0;
  assign reset_values$059 = 5'd0;
  assign reset_values$060 = 5'd0;
  assign reset_values$061 = 5'd0;
  assign reset_values$062 = 5'd0;
  assign reset_values$063 = 5'd0;

  // array declarations
  logic   [   5:0] read_addr[0:0];
  assign read_addr[  0] = read_addr$000;
  logic    [   4:0] read_data[0:0];
  assign read_data$000 = read_data[  0];
  logic    [   4:0] regs[0:63];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  assign regs$002 = regs[  2];
  assign regs$003 = regs[  3];
  assign regs$004 = regs[  4];
  assign regs$005 = regs[  5];
  assign regs$006 = regs[  6];
  assign regs$007 = regs[  7];
  assign regs$008 = regs[  8];
  assign regs$009 = regs[  9];
  assign regs$010 = regs[ 10];
  assign regs$011 = regs[ 11];
  assign regs$012 = regs[ 12];
  assign regs$013 = regs[ 13];
  assign regs$014 = regs[ 14];
  assign regs$015 = regs[ 15];
  assign regs$016 = regs[ 16];
  assign regs$017 = regs[ 17];
  assign regs$018 = regs[ 18];
  assign regs$019 = regs[ 19];
  assign regs$020 = regs[ 20];
  assign regs$021 = regs[ 21];
  assign regs$022 = regs[ 22];
  assign regs$023 = regs[ 23];
  assign regs$024 = regs[ 24];
  assign regs$025 = regs[ 25];
  assign regs$026 = regs[ 26];
  assign regs$027 = regs[ 27];
  assign regs$028 = regs[ 28];
  assign regs$029 = regs[ 29];
  assign regs$030 = regs[ 30];
  assign regs$031 = regs[ 31];
  assign regs$032 = regs[ 32];
  assign regs$033 = regs[ 33];
  assign regs$034 = regs[ 34];
  assign regs$035 = regs[ 35];
  assign regs$036 = regs[ 36];
  assign regs$037 = regs[ 37];
  assign regs$038 = regs[ 38];
  assign regs$039 = regs[ 39];
  assign regs$040 = regs[ 40];
  assign regs$041 = regs[ 41];
  assign regs$042 = regs[ 42];
  assign regs$043 = regs[ 43];
  assign regs$044 = regs[ 44];
  assign regs$045 = regs[ 45];
  assign regs$046 = regs[ 46];
  assign regs$047 = regs[ 47];
  assign regs$048 = regs[ 48];
  assign regs$049 = regs[ 49];
  assign regs$050 = regs[ 50];
  assign regs$051 = regs[ 51];
  assign regs$052 = regs[ 52];
  assign regs$053 = regs[ 53];
  assign regs$054 = regs[ 54];
  assign regs$055 = regs[ 55];
  assign regs$056 = regs[ 56];
  assign regs$057 = regs[ 57];
  assign regs$058 = regs[ 58];
  assign regs$059 = regs[ 59];
  assign regs$060 = regs[ 60];
  assign regs$061 = regs[ 61];
  assign regs$062 = regs[ 62];
  assign regs$063 = regs[ 63];
  logic   [   4:0] reset_values[0:63];
  assign reset_values[  0] = reset_values$000;
  assign reset_values[  1] = reset_values$001;
  assign reset_values[  2] = reset_values$002;
  assign reset_values[  3] = reset_values$003;
  assign reset_values[  4] = reset_values$004;
  assign reset_values[  5] = reset_values$005;
  assign reset_values[  6] = reset_values$006;
  assign reset_values[  7] = reset_values$007;
  assign reset_values[  8] = reset_values$008;
  assign reset_values[  9] = reset_values$009;
  assign reset_values[ 10] = reset_values$010;
  assign reset_values[ 11] = reset_values$011;
  assign reset_values[ 12] = reset_values$012;
  assign reset_values[ 13] = reset_values$013;
  assign reset_values[ 14] = reset_values$014;
  assign reset_values[ 15] = reset_values$015;
  assign reset_values[ 16] = reset_values$016;
  assign reset_values[ 17] = reset_values$017;
  assign reset_values[ 18] = reset_values$018;
  assign reset_values[ 19] = reset_values$019;
  assign reset_values[ 20] = reset_values$020;
  assign reset_values[ 21] = reset_values$021;
  assign reset_values[ 22] = reset_values$022;
  assign reset_values[ 23] = reset_values$023;
  assign reset_values[ 24] = reset_values$024;
  assign reset_values[ 25] = reset_values$025;
  assign reset_values[ 26] = reset_values$026;
  assign reset_values[ 27] = reset_values$027;
  assign reset_values[ 28] = reset_values$028;
  assign reset_values[ 29] = reset_values$029;
  assign reset_values[ 30] = reset_values$030;
  assign reset_values[ 31] = reset_values$031;
  assign reset_values[ 32] = reset_values$032;
  assign reset_values[ 33] = reset_values$033;
  assign reset_values[ 34] = reset_values$034;
  assign reset_values[ 35] = reset_values$035;
  assign reset_values[ 36] = reset_values$036;
  assign reset_values[ 37] = reset_values$037;
  assign reset_values[ 38] = reset_values$038;
  assign reset_values[ 39] = reset_values$039;
  assign reset_values[ 40] = reset_values$040;
  assign reset_values[ 41] = reset_values$041;
  assign reset_values[ 42] = reset_values$042;
  assign reset_values[ 43] = reset_values$043;
  assign reset_values[ 44] = reset_values$044;
  assign reset_values[ 45] = reset_values$045;
  assign reset_values[ 46] = reset_values$046;
  assign reset_values[ 47] = reset_values$047;
  assign reset_values[ 48] = reset_values$048;
  assign reset_values[ 49] = reset_values$049;
  assign reset_values[ 50] = reset_values$050;
  assign reset_values[ 51] = reset_values$051;
  assign reset_values[ 52] = reset_values$052;
  assign reset_values[ 53] = reset_values$053;
  assign reset_values[ 54] = reset_values$054;
  assign reset_values[ 55] = reset_values$055;
  assign reset_values[ 56] = reset_values$056;
  assign reset_values[ 57] = reset_values$057;
  assign reset_values[ 58] = reset_values$058;
  assign reset_values[ 59] = reset_values$059;
  assign reset_values[ 60] = reset_values$060;
  assign reset_values[ 61] = reset_values$061;
  assign reset_values[ 62] = reset_values$062;
  assign reset_values[ 63] = reset_values$063;
  logic   [   5:0] write_addr[0:0];
  assign write_addr[  0] = write_addr$000;
  logic   [   0:0] write_call[0:0];
  assign write_call[  0] = write_call$000;
  logic   [   4:0] write_data[0:0];
  assign write_data[  0] = write_data$000;

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def handle_writes():
  //         if s.reset:
  //           for i in range(nwords):
  //             s.regs[i].n = s.reset_values[i]
  //         else:
  //           for i in range(num_write_ports):
  //             if s.write_call[i]:
  //               s.regs[s.write_addr[i]].n = s.write_data[i]

  // logic for handle_writes()
  always @ (posedge clk) begin
    if (reset) begin
      for (i=0; i < nwords; i=i+1)
      begin
        regs[i] <= reset_values[i];
      end
    end
    else begin
      for (i=0; i < num_write_ports; i=i+1)
      begin
        if (write_call[i]) begin
          regs[write_addr[i]] <= write_data[i];
        end
        else begin
        end
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_reads():
  //         for i in range(num_read_ports):
  //           s.read_data[i].v = s.regs[s.read_addr[i]]
  //           # Bypass logic
  //           for j in range(num_write_ports):
  //             if s.write_call[j] and s.write_addr[j] == s.read_addr[i]:
  //               s.read_data[i].v = s.write_data[j]

  // logic for handle_reads()
  always @ (*) begin
    for (i=0; i < num_read_ports; i=i+1)
    begin
      read_data[i] = regs[read_addr[i]];
      for (j=0; j < num_write_ports; j=j+1)
      begin
        if ((write_call[j]&&(write_addr[j] == read_addr[i]))) begin
          read_data[i] = write_data[j];
        end
        else begin
        end
      end
    end
  end


endmodule // AsynchronousRAM_0x6ff7d20a35694d13

//-----------------------------------------------------------------------------
// RegisterFile_0x6ba986f42995f7d7
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.registerfile {"dtype": 6, "nregs": 32, "num_read_ports": 1, "num_write_ports": 1, "reset_values": [0, 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30], "write_dump_bypass": true, "write_read_bypass": false}
// PyMTL: verilator_xinit = zeros
module RegisterFile_0x6ba986f42995f7d7
(
  input  logic [   0:0] clk,
  output logic [   5:0] dump_out$000,
  output logic [   5:0] dump_out$010,
  output logic [   5:0] dump_out$011,
  output logic [   5:0] dump_out$012,
  output logic [   5:0] dump_out$013,
  output logic [   5:0] dump_out$014,
  output logic [   5:0] dump_out$015,
  output logic [   5:0] dump_out$016,
  output logic [   5:0] dump_out$017,
  output logic [   5:0] dump_out$018,
  output logic [   5:0] dump_out$019,
  output logic [   5:0] dump_out$001,
  output logic [   5:0] dump_out$020,
  output logic [   5:0] dump_out$021,
  output logic [   5:0] dump_out$022,
  output logic [   5:0] dump_out$023,
  output logic [   5:0] dump_out$024,
  output logic [   5:0] dump_out$025,
  output logic [   5:0] dump_out$026,
  output logic [   5:0] dump_out$027,
  output logic [   5:0] dump_out$028,
  output logic [   5:0] dump_out$029,
  output logic [   5:0] dump_out$002,
  output logic [   5:0] dump_out$030,
  output logic [   5:0] dump_out$031,
  output logic [   5:0] dump_out$003,
  output logic [   5:0] dump_out$004,
  output logic [   5:0] dump_out$005,
  output logic [   5:0] dump_out$006,
  output logic [   5:0] dump_out$007,
  output logic [   5:0] dump_out$008,
  output logic [   5:0] dump_out$009,
  input  logic [   4:0] read_addr$000,
  output logic [   5:0] read_data$000,
  input  logic [   0:0] reset,
  input  logic [   0:0] set_call,
  input  logic [   5:0] set_in_$000,
  input  logic [   5:0] set_in_$010,
  input  logic [   5:0] set_in_$011,
  input  logic [   5:0] set_in_$012,
  input  logic [   5:0] set_in_$013,
  input  logic [   5:0] set_in_$014,
  input  logic [   5:0] set_in_$015,
  input  logic [   5:0] set_in_$016,
  input  logic [   5:0] set_in_$017,
  input  logic [   5:0] set_in_$018,
  input  logic [   5:0] set_in_$019,
  input  logic [   5:0] set_in_$001,
  input  logic [   5:0] set_in_$020,
  input  logic [   5:0] set_in_$021,
  input  logic [   5:0] set_in_$022,
  input  logic [   5:0] set_in_$023,
  input  logic [   5:0] set_in_$024,
  input  logic [   5:0] set_in_$025,
  input  logic [   5:0] set_in_$026,
  input  logic [   5:0] set_in_$027,
  input  logic [   5:0] set_in_$028,
  input  logic [   5:0] set_in_$029,
  input  logic [   5:0] set_in_$002,
  input  logic [   5:0] set_in_$030,
  input  logic [   5:0] set_in_$031,
  input  logic [   5:0] set_in_$003,
  input  logic [   5:0] set_in_$004,
  input  logic [   5:0] set_in_$005,
  input  logic [   5:0] set_in_$006,
  input  logic [   5:0] set_in_$007,
  input  logic [   5:0] set_in_$008,
  input  logic [   5:0] set_in_$009,
  input  logic [   4:0] write_addr$000,
  input  logic [   0:0] write_call$000,
  input  logic [   5:0] write_data$000
);

  // logic declarations
  logic   [   5:0] write_inc$000;
  logic   [   5:0] write_inc$001;
  logic   [   5:0] write_inc$002;
  logic   [   5:0] write_inc$003;
  logic   [   5:0] write_inc$004;
  logic   [   5:0] write_inc$005;
  logic   [   5:0] write_inc$006;
  logic   [   5:0] write_inc$007;
  logic   [   5:0] write_inc$008;
  logic   [   5:0] write_inc$009;
  logic   [   5:0] write_inc$010;
  logic   [   5:0] write_inc$011;
  logic   [   5:0] write_inc$012;
  logic   [   5:0] write_inc$013;
  logic   [   5:0] write_inc$014;
  logic   [   5:0] write_inc$015;
  logic   [   5:0] write_inc$016;
  logic   [   5:0] write_inc$017;
  logic   [   5:0] write_inc$018;
  logic   [   5:0] write_inc$019;
  logic   [   5:0] write_inc$020;
  logic   [   5:0] write_inc$021;
  logic   [   5:0] write_inc$022;
  logic   [   5:0] write_inc$023;
  logic   [   5:0] write_inc$024;
  logic   [   5:0] write_inc$025;
  logic   [   5:0] write_inc$026;
  logic   [   5:0] write_inc$027;
  logic   [   5:0] write_inc$028;
  logic   [   5:0] write_inc$029;
  logic   [   5:0] write_inc$030;
  logic   [   5:0] write_inc$031;
  logic   [   5:0] after_set$000;
  logic   [   5:0] after_set$001;
  logic   [   5:0] after_set$002;
  logic   [   5:0] after_set$003;
  logic   [   5:0] after_set$004;
  logic   [   5:0] after_set$005;
  logic   [   5:0] after_set$006;
  logic   [   5:0] after_set$007;
  logic   [   5:0] after_set$008;
  logic   [   5:0] after_set$009;
  logic   [   5:0] after_set$010;
  logic   [   5:0] after_set$011;
  logic   [   5:0] after_set$012;
  logic   [   5:0] after_set$013;
  logic   [   5:0] after_set$014;
  logic   [   5:0] after_set$015;
  logic   [   5:0] after_set$016;
  logic   [   5:0] after_set$017;
  logic   [   5:0] after_set$018;
  logic   [   5:0] after_set$019;
  logic   [   5:0] after_set$020;
  logic   [   5:0] after_set$021;
  logic   [   5:0] after_set$022;
  logic   [   5:0] after_set$023;
  logic   [   5:0] after_set$024;
  logic   [   5:0] after_set$025;
  logic   [   5:0] after_set$026;
  logic   [   5:0] after_set$027;
  logic   [   5:0] after_set$028;
  logic   [   5:0] after_set$029;
  logic   [   5:0] after_set$030;
  logic   [   5:0] after_set$031;
  logic   [   5:0] regs$000;
  logic   [   5:0] regs$001;
  logic   [   5:0] regs$002;
  logic   [   5:0] regs$003;
  logic   [   5:0] regs$004;
  logic   [   5:0] regs$005;
  logic   [   5:0] regs$006;
  logic   [   5:0] regs$007;
  logic   [   5:0] regs$008;
  logic   [   5:0] regs$009;
  logic   [   5:0] regs$010;
  logic   [   5:0] regs$011;
  logic   [   5:0] regs$012;
  logic   [   5:0] regs$013;
  logic   [   5:0] regs$014;
  logic   [   5:0] regs$015;
  logic   [   5:0] regs$016;
  logic   [   5:0] regs$017;
  logic   [   5:0] regs$018;
  logic   [   5:0] regs$019;
  logic   [   5:0] regs$020;
  logic   [   5:0] regs$021;
  logic   [   5:0] regs$022;
  logic   [   5:0] regs$023;
  logic   [   5:0] regs$024;
  logic   [   5:0] regs$025;
  logic   [   5:0] regs$026;
  logic   [   5:0] regs$027;
  logic   [   5:0] regs$028;
  logic   [   5:0] regs$029;
  logic   [   5:0] regs$030;
  logic   [   5:0] regs$031;
  logic   [   5:0] after_write$000;
  logic   [   5:0] after_write$001;
  logic   [   5:0] after_write$002;
  logic   [   5:0] after_write$003;
  logic   [   5:0] after_write$004;
  logic   [   5:0] after_write$005;
  logic   [   5:0] after_write$006;
  logic   [   5:0] after_write$007;
  logic   [   5:0] after_write$008;
  logic   [   5:0] after_write$009;
  logic   [   5:0] after_write$010;
  logic   [   5:0] after_write$011;
  logic   [   5:0] after_write$012;
  logic   [   5:0] after_write$013;
  logic   [   5:0] after_write$014;
  logic   [   5:0] after_write$015;
  logic   [   5:0] after_write$016;
  logic   [   5:0] after_write$017;
  logic   [   5:0] after_write$018;
  logic   [   5:0] after_write$019;
  logic   [   5:0] after_write$020;
  logic   [   5:0] after_write$021;
  logic   [   5:0] after_write$022;
  logic   [   5:0] after_write$023;
  logic   [   5:0] after_write$024;
  logic   [   5:0] after_write$025;
  logic   [   5:0] after_write$026;
  logic   [   5:0] after_write$027;
  logic   [   5:0] after_write$028;
  logic   [   5:0] after_write$029;
  logic   [   5:0] after_write$030;
  logic   [   5:0] after_write$031;


  // signal connections
  assign dump_out$000 = after_write$000;
  assign dump_out$001 = after_write$001;
  assign dump_out$002 = after_write$002;
  assign dump_out$003 = after_write$003;
  assign dump_out$004 = after_write$004;
  assign dump_out$005 = after_write$005;
  assign dump_out$006 = after_write$006;
  assign dump_out$007 = after_write$007;
  assign dump_out$008 = after_write$008;
  assign dump_out$009 = after_write$009;
  assign dump_out$010 = after_write$010;
  assign dump_out$011 = after_write$011;
  assign dump_out$012 = after_write$012;
  assign dump_out$013 = after_write$013;
  assign dump_out$014 = after_write$014;
  assign dump_out$015 = after_write$015;
  assign dump_out$016 = after_write$016;
  assign dump_out$017 = after_write$017;
  assign dump_out$018 = after_write$018;
  assign dump_out$019 = after_write$019;
  assign dump_out$020 = after_write$020;
  assign dump_out$021 = after_write$021;
  assign dump_out$022 = after_write$022;
  assign dump_out$023 = after_write$023;
  assign dump_out$024 = after_write$024;
  assign dump_out$025 = after_write$025;
  assign dump_out$026 = after_write$026;
  assign dump_out$027 = after_write$027;
  assign dump_out$028 = after_write$028;
  assign dump_out$029 = after_write$029;
  assign dump_out$030 = after_write$030;
  assign dump_out$031 = after_write$031;

  // array declarations
  logic    [   5:0] after_set[0:31];
  assign after_set$000 = after_set[  0];
  assign after_set$001 = after_set[  1];
  assign after_set$002 = after_set[  2];
  assign after_set$003 = after_set[  3];
  assign after_set$004 = after_set[  4];
  assign after_set$005 = after_set[  5];
  assign after_set$006 = after_set[  6];
  assign after_set$007 = after_set[  7];
  assign after_set$008 = after_set[  8];
  assign after_set$009 = after_set[  9];
  assign after_set$010 = after_set[ 10];
  assign after_set$011 = after_set[ 11];
  assign after_set$012 = after_set[ 12];
  assign after_set$013 = after_set[ 13];
  assign after_set$014 = after_set[ 14];
  assign after_set$015 = after_set[ 15];
  assign after_set$016 = after_set[ 16];
  assign after_set$017 = after_set[ 17];
  assign after_set$018 = after_set[ 18];
  assign after_set$019 = after_set[ 19];
  assign after_set$020 = after_set[ 20];
  assign after_set$021 = after_set[ 21];
  assign after_set$022 = after_set[ 22];
  assign after_set$023 = after_set[ 23];
  assign after_set$024 = after_set[ 24];
  assign after_set$025 = after_set[ 25];
  assign after_set$026 = after_set[ 26];
  assign after_set$027 = after_set[ 27];
  assign after_set$028 = after_set[ 28];
  assign after_set$029 = after_set[ 29];
  assign after_set$030 = after_set[ 30];
  assign after_set$031 = after_set[ 31];
  logic    [   5:0] after_write[0:31];
  assign after_write$000 = after_write[  0];
  assign after_write$001 = after_write[  1];
  assign after_write$002 = after_write[  2];
  assign after_write$003 = after_write[  3];
  assign after_write$004 = after_write[  4];
  assign after_write$005 = after_write[  5];
  assign after_write$006 = after_write[  6];
  assign after_write$007 = after_write[  7];
  assign after_write$008 = after_write[  8];
  assign after_write$009 = after_write[  9];
  assign after_write$010 = after_write[ 10];
  assign after_write$011 = after_write[ 11];
  assign after_write$012 = after_write[ 12];
  assign after_write$013 = after_write[ 13];
  assign after_write$014 = after_write[ 14];
  assign after_write$015 = after_write[ 15];
  assign after_write$016 = after_write[ 16];
  assign after_write$017 = after_write[ 17];
  assign after_write$018 = after_write[ 18];
  assign after_write$019 = after_write[ 19];
  assign after_write$020 = after_write[ 20];
  assign after_write$021 = after_write[ 21];
  assign after_write$022 = after_write[ 22];
  assign after_write$023 = after_write[ 23];
  assign after_write$024 = after_write[ 24];
  assign after_write$025 = after_write[ 25];
  assign after_write$026 = after_write[ 26];
  assign after_write$027 = after_write[ 27];
  assign after_write$028 = after_write[ 28];
  assign after_write$029 = after_write[ 29];
  assign after_write$030 = after_write[ 30];
  assign after_write$031 = after_write[ 31];
  logic   [   4:0] read_addr[0:0];
  assign read_addr[  0] = read_addr$000;
  logic    [   5:0] read_data[0:0];
  assign read_data$000 = read_data[  0];
  logic    [   5:0] regs[0:31];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  assign regs$002 = regs[  2];
  assign regs$003 = regs[  3];
  assign regs$004 = regs[  4];
  assign regs$005 = regs[  5];
  assign regs$006 = regs[  6];
  assign regs$007 = regs[  7];
  assign regs$008 = regs[  8];
  assign regs$009 = regs[  9];
  assign regs$010 = regs[ 10];
  assign regs$011 = regs[ 11];
  assign regs$012 = regs[ 12];
  assign regs$013 = regs[ 13];
  assign regs$014 = regs[ 14];
  assign regs$015 = regs[ 15];
  assign regs$016 = regs[ 16];
  assign regs$017 = regs[ 17];
  assign regs$018 = regs[ 18];
  assign regs$019 = regs[ 19];
  assign regs$020 = regs[ 20];
  assign regs$021 = regs[ 21];
  assign regs$022 = regs[ 22];
  assign regs$023 = regs[ 23];
  assign regs$024 = regs[ 24];
  assign regs$025 = regs[ 25];
  assign regs$026 = regs[ 26];
  assign regs$027 = regs[ 27];
  assign regs$028 = regs[ 28];
  assign regs$029 = regs[ 29];
  assign regs$030 = regs[ 30];
  assign regs$031 = regs[ 31];
  logic   [   5:0] set_in_[0:31];
  assign set_in_[  0] = set_in_$000;
  assign set_in_[  1] = set_in_$001;
  assign set_in_[  2] = set_in_$002;
  assign set_in_[  3] = set_in_$003;
  assign set_in_[  4] = set_in_$004;
  assign set_in_[  5] = set_in_$005;
  assign set_in_[  6] = set_in_$006;
  assign set_in_[  7] = set_in_$007;
  assign set_in_[  8] = set_in_$008;
  assign set_in_[  9] = set_in_$009;
  assign set_in_[ 10] = set_in_$010;
  assign set_in_[ 11] = set_in_$011;
  assign set_in_[ 12] = set_in_$012;
  assign set_in_[ 13] = set_in_$013;
  assign set_in_[ 14] = set_in_$014;
  assign set_in_[ 15] = set_in_$015;
  assign set_in_[ 16] = set_in_$016;
  assign set_in_[ 17] = set_in_$017;
  assign set_in_[ 18] = set_in_$018;
  assign set_in_[ 19] = set_in_$019;
  assign set_in_[ 20] = set_in_$020;
  assign set_in_[ 21] = set_in_$021;
  assign set_in_[ 22] = set_in_$022;
  assign set_in_[ 23] = set_in_$023;
  assign set_in_[ 24] = set_in_$024;
  assign set_in_[ 25] = set_in_$025;
  assign set_in_[ 26] = set_in_$026;
  assign set_in_[ 27] = set_in_$027;
  assign set_in_[ 28] = set_in_$028;
  assign set_in_[ 29] = set_in_$029;
  assign set_in_[ 30] = set_in_$030;
  assign set_in_[ 31] = set_in_$031;
  logic   [   4:0] write_addr[0:0];
  assign write_addr[  0] = write_addr$000;
  logic   [   0:0] write_call[0:0];
  assign write_call[  0] = write_call$000;
  logic   [   5:0] write_data[0:0];
  assign write_data[  0] = write_data$000;
  logic    [   5:0] write_inc[0:31];
  assign write_inc$000 = write_inc[  0];
  assign write_inc$001 = write_inc[  1];
  assign write_inc$002 = write_inc[  2];
  assign write_inc$003 = write_inc[  3];
  assign write_inc$004 = write_inc[  4];
  assign write_inc$005 = write_inc[  5];
  assign write_inc$006 = write_inc[  6];
  assign write_inc$007 = write_inc[  7];
  assign write_inc$008 = write_inc[  8];
  assign write_inc$009 = write_inc[  9];
  assign write_inc$010 = write_inc[ 10];
  assign write_inc$011 = write_inc[ 11];
  assign write_inc$012 = write_inc[ 12];
  assign write_inc$013 = write_inc[ 13];
  assign write_inc$014 = write_inc[ 14];
  assign write_inc$015 = write_inc[ 15];
  assign write_inc$016 = write_inc[ 16];
  assign write_inc$017 = write_inc[ 17];
  assign write_inc$018 = write_inc[ 18];
  assign write_inc$019 = write_inc[ 19];
  assign write_inc$020 = write_inc[ 20];
  assign write_inc$021 = write_inc[ 21];
  assign write_inc$022 = write_inc[ 22];
  assign write_inc$023 = write_inc[ 23];
  assign write_inc$024 = write_inc[ 24];
  assign write_inc$025 = write_inc[ 25];
  assign write_inc$026 = write_inc[ 26];
  assign write_inc$027 = write_inc[ 27];
  assign write_inc$028 = write_inc[ 28];
  assign write_inc$029 = write_inc[ 29];
  assign write_inc$030 = write_inc[ 30];
  assign write_inc$031 = write_inc[ 31];

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[0] <= 0;
    end
    else begin
      regs[0] <= after_set[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[1] <= 0;
    end
    else begin
      regs[1] <= after_set[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[2] <= 1;
    end
    else begin
      regs[2] <= after_set[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[3] <= 2;
    end
    else begin
      regs[3] <= after_set[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[4] <= 3;
    end
    else begin
      regs[4] <= after_set[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[5] <= 4;
    end
    else begin
      regs[5] <= after_set[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[6] <= 5;
    end
    else begin
      regs[6] <= after_set[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[7] <= 6;
    end
    else begin
      regs[7] <= after_set[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[8] <= 7;
    end
    else begin
      regs[8] <= after_set[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[9] <= 8;
    end
    else begin
      regs[9] <= after_set[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[10] <= 9;
    end
    else begin
      regs[10] <= after_set[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[11] <= 10;
    end
    else begin
      regs[11] <= after_set[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[12] <= 11;
    end
    else begin
      regs[12] <= after_set[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[13] <= 12;
    end
    else begin
      regs[13] <= after_set[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[14] <= 13;
    end
    else begin
      regs[14] <= after_set[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[15] <= 14;
    end
    else begin
      regs[15] <= after_set[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[16] <= 15;
    end
    else begin
      regs[16] <= after_set[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[17] <= 16;
    end
    else begin
      regs[17] <= after_set[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[18] <= 17;
    end
    else begin
      regs[18] <= after_set[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[19] <= 18;
    end
    else begin
      regs[19] <= after_set[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[20] <= 19;
    end
    else begin
      regs[20] <= after_set[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[21] <= 20;
    end
    else begin
      regs[21] <= after_set[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[22] <= 21;
    end
    else begin
      regs[22] <= after_set[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[23] <= 22;
    end
    else begin
      regs[23] <= after_set[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[24] <= 23;
    end
    else begin
      regs[24] <= after_set[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[25] <= 24;
    end
    else begin
      regs[25] <= after_set[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[26] <= 25;
    end
    else begin
      regs[26] <= after_set[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[27] <= 26;
    end
    else begin
      regs[27] <= after_set[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[28] <= 27;
    end
    else begin
      regs[28] <= after_set[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[29] <= 28;
    end
    else begin
      regs[29] <= after_set[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[30] <= 29;
    end
    else begin
      regs[30] <= after_set[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[31] <= 30;
    end
    else begin
      regs[31] <= after_set[31];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 0))) begin
      write_inc[0] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[0] = regs[0];
      end
      else begin
        write_inc[0] = write_inc[-32];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[0] = write_inc[0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[0] = set_in_[0];
    end
    else begin
      after_set[0] = after_write[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 1))) begin
      write_inc[1] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[1] = regs[1];
      end
      else begin
        write_inc[1] = write_inc[-31];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[1] = write_inc[1];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[1] = set_in_[1];
    end
    else begin
      after_set[1] = after_write[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 2))) begin
      write_inc[2] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[2] = regs[2];
      end
      else begin
        write_inc[2] = write_inc[-30];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[2] = write_inc[2];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[2] = set_in_[2];
    end
    else begin
      after_set[2] = after_write[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 3))) begin
      write_inc[3] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[3] = regs[3];
      end
      else begin
        write_inc[3] = write_inc[-29];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[3] = write_inc[3];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[3] = set_in_[3];
    end
    else begin
      after_set[3] = after_write[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 4))) begin
      write_inc[4] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[4] = regs[4];
      end
      else begin
        write_inc[4] = write_inc[-28];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[4] = write_inc[4];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[4] = set_in_[4];
    end
    else begin
      after_set[4] = after_write[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 5))) begin
      write_inc[5] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[5] = regs[5];
      end
      else begin
        write_inc[5] = write_inc[-27];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[5] = write_inc[5];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[5] = set_in_[5];
    end
    else begin
      after_set[5] = after_write[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 6))) begin
      write_inc[6] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[6] = regs[6];
      end
      else begin
        write_inc[6] = write_inc[-26];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[6] = write_inc[6];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[6] = set_in_[6];
    end
    else begin
      after_set[6] = after_write[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 7))) begin
      write_inc[7] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[7] = regs[7];
      end
      else begin
        write_inc[7] = write_inc[-25];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[7] = write_inc[7];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[7] = set_in_[7];
    end
    else begin
      after_set[7] = after_write[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 8))) begin
      write_inc[8] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[8] = regs[8];
      end
      else begin
        write_inc[8] = write_inc[-24];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[8] = write_inc[8];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[8] = set_in_[8];
    end
    else begin
      after_set[8] = after_write[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 9))) begin
      write_inc[9] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[9] = regs[9];
      end
      else begin
        write_inc[9] = write_inc[-23];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[9] = write_inc[9];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[9] = set_in_[9];
    end
    else begin
      after_set[9] = after_write[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 10))) begin
      write_inc[10] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[10] = regs[10];
      end
      else begin
        write_inc[10] = write_inc[-22];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[10] = write_inc[10];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[10] = set_in_[10];
    end
    else begin
      after_set[10] = after_write[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 11))) begin
      write_inc[11] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[11] = regs[11];
      end
      else begin
        write_inc[11] = write_inc[-21];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[11] = write_inc[11];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[11] = set_in_[11];
    end
    else begin
      after_set[11] = after_write[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 12))) begin
      write_inc[12] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[12] = regs[12];
      end
      else begin
        write_inc[12] = write_inc[-20];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[12] = write_inc[12];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[12] = set_in_[12];
    end
    else begin
      after_set[12] = after_write[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 13))) begin
      write_inc[13] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[13] = regs[13];
      end
      else begin
        write_inc[13] = write_inc[-19];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[13] = write_inc[13];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[13] = set_in_[13];
    end
    else begin
      after_set[13] = after_write[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 14))) begin
      write_inc[14] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[14] = regs[14];
      end
      else begin
        write_inc[14] = write_inc[-18];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[14] = write_inc[14];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[14] = set_in_[14];
    end
    else begin
      after_set[14] = after_write[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 15))) begin
      write_inc[15] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[15] = regs[15];
      end
      else begin
        write_inc[15] = write_inc[-17];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[15] = write_inc[15];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[15] = set_in_[15];
    end
    else begin
      after_set[15] = after_write[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 16))) begin
      write_inc[16] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[16] = regs[16];
      end
      else begin
        write_inc[16] = write_inc[-16];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[16] = write_inc[16];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[16] = set_in_[16];
    end
    else begin
      after_set[16] = after_write[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 17))) begin
      write_inc[17] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[17] = regs[17];
      end
      else begin
        write_inc[17] = write_inc[-15];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[17] = write_inc[17];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[17] = set_in_[17];
    end
    else begin
      after_set[17] = after_write[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 18))) begin
      write_inc[18] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[18] = regs[18];
      end
      else begin
        write_inc[18] = write_inc[-14];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[18] = write_inc[18];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[18] = set_in_[18];
    end
    else begin
      after_set[18] = after_write[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 19))) begin
      write_inc[19] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[19] = regs[19];
      end
      else begin
        write_inc[19] = write_inc[-13];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[19] = write_inc[19];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[19] = set_in_[19];
    end
    else begin
      after_set[19] = after_write[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 20))) begin
      write_inc[20] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[20] = regs[20];
      end
      else begin
        write_inc[20] = write_inc[-12];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[20] = write_inc[20];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[20] = set_in_[20];
    end
    else begin
      after_set[20] = after_write[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 21))) begin
      write_inc[21] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[21] = regs[21];
      end
      else begin
        write_inc[21] = write_inc[-11];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[21] = write_inc[21];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[21] = set_in_[21];
    end
    else begin
      after_set[21] = after_write[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 22))) begin
      write_inc[22] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[22] = regs[22];
      end
      else begin
        write_inc[22] = write_inc[-10];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[22] = write_inc[22];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[22] = set_in_[22];
    end
    else begin
      after_set[22] = after_write[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 23))) begin
      write_inc[23] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[23] = regs[23];
      end
      else begin
        write_inc[23] = write_inc[-9];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[23] = write_inc[23];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[23] = set_in_[23];
    end
    else begin
      after_set[23] = after_write[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 24))) begin
      write_inc[24] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[24] = regs[24];
      end
      else begin
        write_inc[24] = write_inc[-8];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[24] = write_inc[24];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[24] = set_in_[24];
    end
    else begin
      after_set[24] = after_write[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 25))) begin
      write_inc[25] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[25] = regs[25];
      end
      else begin
        write_inc[25] = write_inc[-7];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[25] = write_inc[25];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[25] = set_in_[25];
    end
    else begin
      after_set[25] = after_write[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 26))) begin
      write_inc[26] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[26] = regs[26];
      end
      else begin
        write_inc[26] = write_inc[-6];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[26] = write_inc[26];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[26] = set_in_[26];
    end
    else begin
      after_set[26] = after_write[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 27))) begin
      write_inc[27] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[27] = regs[27];
      end
      else begin
        write_inc[27] = write_inc[-5];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[27] = write_inc[27];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[27] = set_in_[27];
    end
    else begin
      after_set[27] = after_write[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 28))) begin
      write_inc[28] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[28] = regs[28];
      end
      else begin
        write_inc[28] = write_inc[-4];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[28] = write_inc[28];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[28] = set_in_[28];
    end
    else begin
      after_set[28] = after_write[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 29))) begin
      write_inc[29] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[29] = regs[29];
      end
      else begin
        write_inc[29] = write_inc[-3];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[29] = write_inc[29];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[29] = set_in_[29];
    end
    else begin
      after_set[29] = after_write[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 30))) begin
      write_inc[30] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[30] = regs[30];
      end
      else begin
        write_inc[30] = write_inc[-2];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[30] = write_inc[30];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[30] = set_in_[30];
    end
    else begin
      after_set[30] = after_write[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 31))) begin
      write_inc[31] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[31] = regs[31];
      end
      else begin
        write_inc[31] = write_inc[-1];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[31] = write_inc[31];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[31] = set_in_[31];
    end
    else begin
      after_set[31] = after_write[31];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_read(port=port):
  //           s.read_data[port].v = s.regs[s.read_addr[port]]

  // logic for handle_read()
  always @ (*) begin
    read_data[0] = regs[read_addr[0]];
  end


endmodule // RegisterFile_0x6ba986f42995f7d7

//-----------------------------------------------------------------------------
// RegisterFile_0x39d647b3aea936a6
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.registerfile {"dtype": 1, "nregs": 63, "num_read_ports": 0, "num_write_ports": 2, "reset_values": ["1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "1", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0", "0"], "write_dump_bypass": true, "write_read_bypass": false}
// PyMTL: verilator_xinit = zeros
module RegisterFile_0x39d647b3aea936a6
(
  input  logic [   0:0] clk,
  output logic [   0:0] dump_out$000,
  output logic [   0:0] dump_out$010,
  output logic [   0:0] dump_out$011,
  output logic [   0:0] dump_out$012,
  output logic [   0:0] dump_out$013,
  output logic [   0:0] dump_out$014,
  output logic [   0:0] dump_out$015,
  output logic [   0:0] dump_out$016,
  output logic [   0:0] dump_out$017,
  output logic [   0:0] dump_out$018,
  output logic [   0:0] dump_out$019,
  output logic [   0:0] dump_out$001,
  output logic [   0:0] dump_out$020,
  output logic [   0:0] dump_out$021,
  output logic [   0:0] dump_out$022,
  output logic [   0:0] dump_out$023,
  output logic [   0:0] dump_out$024,
  output logic [   0:0] dump_out$025,
  output logic [   0:0] dump_out$026,
  output logic [   0:0] dump_out$027,
  output logic [   0:0] dump_out$028,
  output logic [   0:0] dump_out$029,
  output logic [   0:0] dump_out$002,
  output logic [   0:0] dump_out$030,
  output logic [   0:0] dump_out$031,
  output logic [   0:0] dump_out$032,
  output logic [   0:0] dump_out$033,
  output logic [   0:0] dump_out$034,
  output logic [   0:0] dump_out$035,
  output logic [   0:0] dump_out$036,
  output logic [   0:0] dump_out$037,
  output logic [   0:0] dump_out$038,
  output logic [   0:0] dump_out$039,
  output logic [   0:0] dump_out$003,
  output logic [   0:0] dump_out$040,
  output logic [   0:0] dump_out$041,
  output logic [   0:0] dump_out$042,
  output logic [   0:0] dump_out$043,
  output logic [   0:0] dump_out$044,
  output logic [   0:0] dump_out$045,
  output logic [   0:0] dump_out$046,
  output logic [   0:0] dump_out$047,
  output logic [   0:0] dump_out$048,
  output logic [   0:0] dump_out$049,
  output logic [   0:0] dump_out$004,
  output logic [   0:0] dump_out$050,
  output logic [   0:0] dump_out$051,
  output logic [   0:0] dump_out$052,
  output logic [   0:0] dump_out$053,
  output logic [   0:0] dump_out$054,
  output logic [   0:0] dump_out$055,
  output logic [   0:0] dump_out$056,
  output logic [   0:0] dump_out$057,
  output logic [   0:0] dump_out$058,
  output logic [   0:0] dump_out$059,
  output logic [   0:0] dump_out$005,
  output logic [   0:0] dump_out$060,
  output logic [   0:0] dump_out$061,
  output logic [   0:0] dump_out$062,
  output logic [   0:0] dump_out$006,
  output logic [   0:0] dump_out$007,
  output logic [   0:0] dump_out$008,
  output logic [   0:0] dump_out$009,
  input  logic [   0:0] reset,
  input  logic [   0:0] set_call,
  input  logic [   0:0] set_in_$000,
  input  logic [   0:0] set_in_$010,
  input  logic [   0:0] set_in_$011,
  input  logic [   0:0] set_in_$012,
  input  logic [   0:0] set_in_$013,
  input  logic [   0:0] set_in_$014,
  input  logic [   0:0] set_in_$015,
  input  logic [   0:0] set_in_$016,
  input  logic [   0:0] set_in_$017,
  input  logic [   0:0] set_in_$018,
  input  logic [   0:0] set_in_$019,
  input  logic [   0:0] set_in_$001,
  input  logic [   0:0] set_in_$020,
  input  logic [   0:0] set_in_$021,
  input  logic [   0:0] set_in_$022,
  input  logic [   0:0] set_in_$023,
  input  logic [   0:0] set_in_$024,
  input  logic [   0:0] set_in_$025,
  input  logic [   0:0] set_in_$026,
  input  logic [   0:0] set_in_$027,
  input  logic [   0:0] set_in_$028,
  input  logic [   0:0] set_in_$029,
  input  logic [   0:0] set_in_$002,
  input  logic [   0:0] set_in_$030,
  input  logic [   0:0] set_in_$031,
  input  logic [   0:0] set_in_$032,
  input  logic [   0:0] set_in_$033,
  input  logic [   0:0] set_in_$034,
  input  logic [   0:0] set_in_$035,
  input  logic [   0:0] set_in_$036,
  input  logic [   0:0] set_in_$037,
  input  logic [   0:0] set_in_$038,
  input  logic [   0:0] set_in_$039,
  input  logic [   0:0] set_in_$003,
  input  logic [   0:0] set_in_$040,
  input  logic [   0:0] set_in_$041,
  input  logic [   0:0] set_in_$042,
  input  logic [   0:0] set_in_$043,
  input  logic [   0:0] set_in_$044,
  input  logic [   0:0] set_in_$045,
  input  logic [   0:0] set_in_$046,
  input  logic [   0:0] set_in_$047,
  input  logic [   0:0] set_in_$048,
  input  logic [   0:0] set_in_$049,
  input  logic [   0:0] set_in_$004,
  input  logic [   0:0] set_in_$050,
  input  logic [   0:0] set_in_$051,
  input  logic [   0:0] set_in_$052,
  input  logic [   0:0] set_in_$053,
  input  logic [   0:0] set_in_$054,
  input  logic [   0:0] set_in_$055,
  input  logic [   0:0] set_in_$056,
  input  logic [   0:0] set_in_$057,
  input  logic [   0:0] set_in_$058,
  input  logic [   0:0] set_in_$059,
  input  logic [   0:0] set_in_$005,
  input  logic [   0:0] set_in_$060,
  input  logic [   0:0] set_in_$061,
  input  logic [   0:0] set_in_$062,
  input  logic [   0:0] set_in_$006,
  input  logic [   0:0] set_in_$007,
  input  logic [   0:0] set_in_$008,
  input  logic [   0:0] set_in_$009,
  input  logic [   5:0] write_addr$000,
  input  logic [   5:0] write_addr$001,
  input  logic [   0:0] write_call$000,
  input  logic [   0:0] write_call$001,
  input  logic [   0:0] write_data$000,
  input  logic [   0:0] write_data$001
);

  // logic declarations
  logic   [   0:0] write_inc$000;
  logic   [   0:0] write_inc$001;
  logic   [   0:0] write_inc$002;
  logic   [   0:0] write_inc$003;
  logic   [   0:0] write_inc$004;
  logic   [   0:0] write_inc$005;
  logic   [   0:0] write_inc$006;
  logic   [   0:0] write_inc$007;
  logic   [   0:0] write_inc$008;
  logic   [   0:0] write_inc$009;
  logic   [   0:0] write_inc$010;
  logic   [   0:0] write_inc$011;
  logic   [   0:0] write_inc$012;
  logic   [   0:0] write_inc$013;
  logic   [   0:0] write_inc$014;
  logic   [   0:0] write_inc$015;
  logic   [   0:0] write_inc$016;
  logic   [   0:0] write_inc$017;
  logic   [   0:0] write_inc$018;
  logic   [   0:0] write_inc$019;
  logic   [   0:0] write_inc$020;
  logic   [   0:0] write_inc$021;
  logic   [   0:0] write_inc$022;
  logic   [   0:0] write_inc$023;
  logic   [   0:0] write_inc$024;
  logic   [   0:0] write_inc$025;
  logic   [   0:0] write_inc$026;
  logic   [   0:0] write_inc$027;
  logic   [   0:0] write_inc$028;
  logic   [   0:0] write_inc$029;
  logic   [   0:0] write_inc$030;
  logic   [   0:0] write_inc$031;
  logic   [   0:0] write_inc$032;
  logic   [   0:0] write_inc$033;
  logic   [   0:0] write_inc$034;
  logic   [   0:0] write_inc$035;
  logic   [   0:0] write_inc$036;
  logic   [   0:0] write_inc$037;
  logic   [   0:0] write_inc$038;
  logic   [   0:0] write_inc$039;
  logic   [   0:0] write_inc$040;
  logic   [   0:0] write_inc$041;
  logic   [   0:0] write_inc$042;
  logic   [   0:0] write_inc$043;
  logic   [   0:0] write_inc$044;
  logic   [   0:0] write_inc$045;
  logic   [   0:0] write_inc$046;
  logic   [   0:0] write_inc$047;
  logic   [   0:0] write_inc$048;
  logic   [   0:0] write_inc$049;
  logic   [   0:0] write_inc$050;
  logic   [   0:0] write_inc$051;
  logic   [   0:0] write_inc$052;
  logic   [   0:0] write_inc$053;
  logic   [   0:0] write_inc$054;
  logic   [   0:0] write_inc$055;
  logic   [   0:0] write_inc$056;
  logic   [   0:0] write_inc$057;
  logic   [   0:0] write_inc$058;
  logic   [   0:0] write_inc$059;
  logic   [   0:0] write_inc$060;
  logic   [   0:0] write_inc$061;
  logic   [   0:0] write_inc$062;
  logic   [   0:0] write_inc$063;
  logic   [   0:0] write_inc$064;
  logic   [   0:0] write_inc$065;
  logic   [   0:0] write_inc$066;
  logic   [   0:0] write_inc$067;
  logic   [   0:0] write_inc$068;
  logic   [   0:0] write_inc$069;
  logic   [   0:0] write_inc$070;
  logic   [   0:0] write_inc$071;
  logic   [   0:0] write_inc$072;
  logic   [   0:0] write_inc$073;
  logic   [   0:0] write_inc$074;
  logic   [   0:0] write_inc$075;
  logic   [   0:0] write_inc$076;
  logic   [   0:0] write_inc$077;
  logic   [   0:0] write_inc$078;
  logic   [   0:0] write_inc$079;
  logic   [   0:0] write_inc$080;
  logic   [   0:0] write_inc$081;
  logic   [   0:0] write_inc$082;
  logic   [   0:0] write_inc$083;
  logic   [   0:0] write_inc$084;
  logic   [   0:0] write_inc$085;
  logic   [   0:0] write_inc$086;
  logic   [   0:0] write_inc$087;
  logic   [   0:0] write_inc$088;
  logic   [   0:0] write_inc$089;
  logic   [   0:0] write_inc$090;
  logic   [   0:0] write_inc$091;
  logic   [   0:0] write_inc$092;
  logic   [   0:0] write_inc$093;
  logic   [   0:0] write_inc$094;
  logic   [   0:0] write_inc$095;
  logic   [   0:0] write_inc$096;
  logic   [   0:0] write_inc$097;
  logic   [   0:0] write_inc$098;
  logic   [   0:0] write_inc$099;
  logic   [   0:0] write_inc$100;
  logic   [   0:0] write_inc$101;
  logic   [   0:0] write_inc$102;
  logic   [   0:0] write_inc$103;
  logic   [   0:0] write_inc$104;
  logic   [   0:0] write_inc$105;
  logic   [   0:0] write_inc$106;
  logic   [   0:0] write_inc$107;
  logic   [   0:0] write_inc$108;
  logic   [   0:0] write_inc$109;
  logic   [   0:0] write_inc$110;
  logic   [   0:0] write_inc$111;
  logic   [   0:0] write_inc$112;
  logic   [   0:0] write_inc$113;
  logic   [   0:0] write_inc$114;
  logic   [   0:0] write_inc$115;
  logic   [   0:0] write_inc$116;
  logic   [   0:0] write_inc$117;
  logic   [   0:0] write_inc$118;
  logic   [   0:0] write_inc$119;
  logic   [   0:0] write_inc$120;
  logic   [   0:0] write_inc$121;
  logic   [   0:0] write_inc$122;
  logic   [   0:0] write_inc$123;
  logic   [   0:0] write_inc$124;
  logic   [   0:0] write_inc$125;
  logic   [   0:0] after_set$000;
  logic   [   0:0] after_set$001;
  logic   [   0:0] after_set$002;
  logic   [   0:0] after_set$003;
  logic   [   0:0] after_set$004;
  logic   [   0:0] after_set$005;
  logic   [   0:0] after_set$006;
  logic   [   0:0] after_set$007;
  logic   [   0:0] after_set$008;
  logic   [   0:0] after_set$009;
  logic   [   0:0] after_set$010;
  logic   [   0:0] after_set$011;
  logic   [   0:0] after_set$012;
  logic   [   0:0] after_set$013;
  logic   [   0:0] after_set$014;
  logic   [   0:0] after_set$015;
  logic   [   0:0] after_set$016;
  logic   [   0:0] after_set$017;
  logic   [   0:0] after_set$018;
  logic   [   0:0] after_set$019;
  logic   [   0:0] after_set$020;
  logic   [   0:0] after_set$021;
  logic   [   0:0] after_set$022;
  logic   [   0:0] after_set$023;
  logic   [   0:0] after_set$024;
  logic   [   0:0] after_set$025;
  logic   [   0:0] after_set$026;
  logic   [   0:0] after_set$027;
  logic   [   0:0] after_set$028;
  logic   [   0:0] after_set$029;
  logic   [   0:0] after_set$030;
  logic   [   0:0] after_set$031;
  logic   [   0:0] after_set$032;
  logic   [   0:0] after_set$033;
  logic   [   0:0] after_set$034;
  logic   [   0:0] after_set$035;
  logic   [   0:0] after_set$036;
  logic   [   0:0] after_set$037;
  logic   [   0:0] after_set$038;
  logic   [   0:0] after_set$039;
  logic   [   0:0] after_set$040;
  logic   [   0:0] after_set$041;
  logic   [   0:0] after_set$042;
  logic   [   0:0] after_set$043;
  logic   [   0:0] after_set$044;
  logic   [   0:0] after_set$045;
  logic   [   0:0] after_set$046;
  logic   [   0:0] after_set$047;
  logic   [   0:0] after_set$048;
  logic   [   0:0] after_set$049;
  logic   [   0:0] after_set$050;
  logic   [   0:0] after_set$051;
  logic   [   0:0] after_set$052;
  logic   [   0:0] after_set$053;
  logic   [   0:0] after_set$054;
  logic   [   0:0] after_set$055;
  logic   [   0:0] after_set$056;
  logic   [   0:0] after_set$057;
  logic   [   0:0] after_set$058;
  logic   [   0:0] after_set$059;
  logic   [   0:0] after_set$060;
  logic   [   0:0] after_set$061;
  logic   [   0:0] after_set$062;
  logic   [   0:0] regs$000;
  logic   [   0:0] regs$001;
  logic   [   0:0] regs$002;
  logic   [   0:0] regs$003;
  logic   [   0:0] regs$004;
  logic   [   0:0] regs$005;
  logic   [   0:0] regs$006;
  logic   [   0:0] regs$007;
  logic   [   0:0] regs$008;
  logic   [   0:0] regs$009;
  logic   [   0:0] regs$010;
  logic   [   0:0] regs$011;
  logic   [   0:0] regs$012;
  logic   [   0:0] regs$013;
  logic   [   0:0] regs$014;
  logic   [   0:0] regs$015;
  logic   [   0:0] regs$016;
  logic   [   0:0] regs$017;
  logic   [   0:0] regs$018;
  logic   [   0:0] regs$019;
  logic   [   0:0] regs$020;
  logic   [   0:0] regs$021;
  logic   [   0:0] regs$022;
  logic   [   0:0] regs$023;
  logic   [   0:0] regs$024;
  logic   [   0:0] regs$025;
  logic   [   0:0] regs$026;
  logic   [   0:0] regs$027;
  logic   [   0:0] regs$028;
  logic   [   0:0] regs$029;
  logic   [   0:0] regs$030;
  logic   [   0:0] regs$031;
  logic   [   0:0] regs$032;
  logic   [   0:0] regs$033;
  logic   [   0:0] regs$034;
  logic   [   0:0] regs$035;
  logic   [   0:0] regs$036;
  logic   [   0:0] regs$037;
  logic   [   0:0] regs$038;
  logic   [   0:0] regs$039;
  logic   [   0:0] regs$040;
  logic   [   0:0] regs$041;
  logic   [   0:0] regs$042;
  logic   [   0:0] regs$043;
  logic   [   0:0] regs$044;
  logic   [   0:0] regs$045;
  logic   [   0:0] regs$046;
  logic   [   0:0] regs$047;
  logic   [   0:0] regs$048;
  logic   [   0:0] regs$049;
  logic   [   0:0] regs$050;
  logic   [   0:0] regs$051;
  logic   [   0:0] regs$052;
  logic   [   0:0] regs$053;
  logic   [   0:0] regs$054;
  logic   [   0:0] regs$055;
  logic   [   0:0] regs$056;
  logic   [   0:0] regs$057;
  logic   [   0:0] regs$058;
  logic   [   0:0] regs$059;
  logic   [   0:0] regs$060;
  logic   [   0:0] regs$061;
  logic   [   0:0] regs$062;
  logic   [   0:0] after_write$000;
  logic   [   0:0] after_write$001;
  logic   [   0:0] after_write$002;
  logic   [   0:0] after_write$003;
  logic   [   0:0] after_write$004;
  logic   [   0:0] after_write$005;
  logic   [   0:0] after_write$006;
  logic   [   0:0] after_write$007;
  logic   [   0:0] after_write$008;
  logic   [   0:0] after_write$009;
  logic   [   0:0] after_write$010;
  logic   [   0:0] after_write$011;
  logic   [   0:0] after_write$012;
  logic   [   0:0] after_write$013;
  logic   [   0:0] after_write$014;
  logic   [   0:0] after_write$015;
  logic   [   0:0] after_write$016;
  logic   [   0:0] after_write$017;
  logic   [   0:0] after_write$018;
  logic   [   0:0] after_write$019;
  logic   [   0:0] after_write$020;
  logic   [   0:0] after_write$021;
  logic   [   0:0] after_write$022;
  logic   [   0:0] after_write$023;
  logic   [   0:0] after_write$024;
  logic   [   0:0] after_write$025;
  logic   [   0:0] after_write$026;
  logic   [   0:0] after_write$027;
  logic   [   0:0] after_write$028;
  logic   [   0:0] after_write$029;
  logic   [   0:0] after_write$030;
  logic   [   0:0] after_write$031;
  logic   [   0:0] after_write$032;
  logic   [   0:0] after_write$033;
  logic   [   0:0] after_write$034;
  logic   [   0:0] after_write$035;
  logic   [   0:0] after_write$036;
  logic   [   0:0] after_write$037;
  logic   [   0:0] after_write$038;
  logic   [   0:0] after_write$039;
  logic   [   0:0] after_write$040;
  logic   [   0:0] after_write$041;
  logic   [   0:0] after_write$042;
  logic   [   0:0] after_write$043;
  logic   [   0:0] after_write$044;
  logic   [   0:0] after_write$045;
  logic   [   0:0] after_write$046;
  logic   [   0:0] after_write$047;
  logic   [   0:0] after_write$048;
  logic   [   0:0] after_write$049;
  logic   [   0:0] after_write$050;
  logic   [   0:0] after_write$051;
  logic   [   0:0] after_write$052;
  logic   [   0:0] after_write$053;
  logic   [   0:0] after_write$054;
  logic   [   0:0] after_write$055;
  logic   [   0:0] after_write$056;
  logic   [   0:0] after_write$057;
  logic   [   0:0] after_write$058;
  logic   [   0:0] after_write$059;
  logic   [   0:0] after_write$060;
  logic   [   0:0] after_write$061;
  logic   [   0:0] after_write$062;


  // signal connections
  assign dump_out$000 = after_write$000;
  assign dump_out$001 = after_write$001;
  assign dump_out$002 = after_write$002;
  assign dump_out$003 = after_write$003;
  assign dump_out$004 = after_write$004;
  assign dump_out$005 = after_write$005;
  assign dump_out$006 = after_write$006;
  assign dump_out$007 = after_write$007;
  assign dump_out$008 = after_write$008;
  assign dump_out$009 = after_write$009;
  assign dump_out$010 = after_write$010;
  assign dump_out$011 = after_write$011;
  assign dump_out$012 = after_write$012;
  assign dump_out$013 = after_write$013;
  assign dump_out$014 = after_write$014;
  assign dump_out$015 = after_write$015;
  assign dump_out$016 = after_write$016;
  assign dump_out$017 = after_write$017;
  assign dump_out$018 = after_write$018;
  assign dump_out$019 = after_write$019;
  assign dump_out$020 = after_write$020;
  assign dump_out$021 = after_write$021;
  assign dump_out$022 = after_write$022;
  assign dump_out$023 = after_write$023;
  assign dump_out$024 = after_write$024;
  assign dump_out$025 = after_write$025;
  assign dump_out$026 = after_write$026;
  assign dump_out$027 = after_write$027;
  assign dump_out$028 = after_write$028;
  assign dump_out$029 = after_write$029;
  assign dump_out$030 = after_write$030;
  assign dump_out$031 = after_write$031;
  assign dump_out$032 = after_write$032;
  assign dump_out$033 = after_write$033;
  assign dump_out$034 = after_write$034;
  assign dump_out$035 = after_write$035;
  assign dump_out$036 = after_write$036;
  assign dump_out$037 = after_write$037;
  assign dump_out$038 = after_write$038;
  assign dump_out$039 = after_write$039;
  assign dump_out$040 = after_write$040;
  assign dump_out$041 = after_write$041;
  assign dump_out$042 = after_write$042;
  assign dump_out$043 = after_write$043;
  assign dump_out$044 = after_write$044;
  assign dump_out$045 = after_write$045;
  assign dump_out$046 = after_write$046;
  assign dump_out$047 = after_write$047;
  assign dump_out$048 = after_write$048;
  assign dump_out$049 = after_write$049;
  assign dump_out$050 = after_write$050;
  assign dump_out$051 = after_write$051;
  assign dump_out$052 = after_write$052;
  assign dump_out$053 = after_write$053;
  assign dump_out$054 = after_write$054;
  assign dump_out$055 = after_write$055;
  assign dump_out$056 = after_write$056;
  assign dump_out$057 = after_write$057;
  assign dump_out$058 = after_write$058;
  assign dump_out$059 = after_write$059;
  assign dump_out$060 = after_write$060;
  assign dump_out$061 = after_write$061;
  assign dump_out$062 = after_write$062;

  // array declarations
  logic    [   0:0] after_set[0:62];
  assign after_set$000 = after_set[  0];
  assign after_set$001 = after_set[  1];
  assign after_set$002 = after_set[  2];
  assign after_set$003 = after_set[  3];
  assign after_set$004 = after_set[  4];
  assign after_set$005 = after_set[  5];
  assign after_set$006 = after_set[  6];
  assign after_set$007 = after_set[  7];
  assign after_set$008 = after_set[  8];
  assign after_set$009 = after_set[  9];
  assign after_set$010 = after_set[ 10];
  assign after_set$011 = after_set[ 11];
  assign after_set$012 = after_set[ 12];
  assign after_set$013 = after_set[ 13];
  assign after_set$014 = after_set[ 14];
  assign after_set$015 = after_set[ 15];
  assign after_set$016 = after_set[ 16];
  assign after_set$017 = after_set[ 17];
  assign after_set$018 = after_set[ 18];
  assign after_set$019 = after_set[ 19];
  assign after_set$020 = after_set[ 20];
  assign after_set$021 = after_set[ 21];
  assign after_set$022 = after_set[ 22];
  assign after_set$023 = after_set[ 23];
  assign after_set$024 = after_set[ 24];
  assign after_set$025 = after_set[ 25];
  assign after_set$026 = after_set[ 26];
  assign after_set$027 = after_set[ 27];
  assign after_set$028 = after_set[ 28];
  assign after_set$029 = after_set[ 29];
  assign after_set$030 = after_set[ 30];
  assign after_set$031 = after_set[ 31];
  assign after_set$032 = after_set[ 32];
  assign after_set$033 = after_set[ 33];
  assign after_set$034 = after_set[ 34];
  assign after_set$035 = after_set[ 35];
  assign after_set$036 = after_set[ 36];
  assign after_set$037 = after_set[ 37];
  assign after_set$038 = after_set[ 38];
  assign after_set$039 = after_set[ 39];
  assign after_set$040 = after_set[ 40];
  assign after_set$041 = after_set[ 41];
  assign after_set$042 = after_set[ 42];
  assign after_set$043 = after_set[ 43];
  assign after_set$044 = after_set[ 44];
  assign after_set$045 = after_set[ 45];
  assign after_set$046 = after_set[ 46];
  assign after_set$047 = after_set[ 47];
  assign after_set$048 = after_set[ 48];
  assign after_set$049 = after_set[ 49];
  assign after_set$050 = after_set[ 50];
  assign after_set$051 = after_set[ 51];
  assign after_set$052 = after_set[ 52];
  assign after_set$053 = after_set[ 53];
  assign after_set$054 = after_set[ 54];
  assign after_set$055 = after_set[ 55];
  assign after_set$056 = after_set[ 56];
  assign after_set$057 = after_set[ 57];
  assign after_set$058 = after_set[ 58];
  assign after_set$059 = after_set[ 59];
  assign after_set$060 = after_set[ 60];
  assign after_set$061 = after_set[ 61];
  assign after_set$062 = after_set[ 62];
  logic    [   0:0] after_write[0:62];
  assign after_write$000 = after_write[  0];
  assign after_write$001 = after_write[  1];
  assign after_write$002 = after_write[  2];
  assign after_write$003 = after_write[  3];
  assign after_write$004 = after_write[  4];
  assign after_write$005 = after_write[  5];
  assign after_write$006 = after_write[  6];
  assign after_write$007 = after_write[  7];
  assign after_write$008 = after_write[  8];
  assign after_write$009 = after_write[  9];
  assign after_write$010 = after_write[ 10];
  assign after_write$011 = after_write[ 11];
  assign after_write$012 = after_write[ 12];
  assign after_write$013 = after_write[ 13];
  assign after_write$014 = after_write[ 14];
  assign after_write$015 = after_write[ 15];
  assign after_write$016 = after_write[ 16];
  assign after_write$017 = after_write[ 17];
  assign after_write$018 = after_write[ 18];
  assign after_write$019 = after_write[ 19];
  assign after_write$020 = after_write[ 20];
  assign after_write$021 = after_write[ 21];
  assign after_write$022 = after_write[ 22];
  assign after_write$023 = after_write[ 23];
  assign after_write$024 = after_write[ 24];
  assign after_write$025 = after_write[ 25];
  assign after_write$026 = after_write[ 26];
  assign after_write$027 = after_write[ 27];
  assign after_write$028 = after_write[ 28];
  assign after_write$029 = after_write[ 29];
  assign after_write$030 = after_write[ 30];
  assign after_write$031 = after_write[ 31];
  assign after_write$032 = after_write[ 32];
  assign after_write$033 = after_write[ 33];
  assign after_write$034 = after_write[ 34];
  assign after_write$035 = after_write[ 35];
  assign after_write$036 = after_write[ 36];
  assign after_write$037 = after_write[ 37];
  assign after_write$038 = after_write[ 38];
  assign after_write$039 = after_write[ 39];
  assign after_write$040 = after_write[ 40];
  assign after_write$041 = after_write[ 41];
  assign after_write$042 = after_write[ 42];
  assign after_write$043 = after_write[ 43];
  assign after_write$044 = after_write[ 44];
  assign after_write$045 = after_write[ 45];
  assign after_write$046 = after_write[ 46];
  assign after_write$047 = after_write[ 47];
  assign after_write$048 = after_write[ 48];
  assign after_write$049 = after_write[ 49];
  assign after_write$050 = after_write[ 50];
  assign after_write$051 = after_write[ 51];
  assign after_write$052 = after_write[ 52];
  assign after_write$053 = after_write[ 53];
  assign after_write$054 = after_write[ 54];
  assign after_write$055 = after_write[ 55];
  assign after_write$056 = after_write[ 56];
  assign after_write$057 = after_write[ 57];
  assign after_write$058 = after_write[ 58];
  assign after_write$059 = after_write[ 59];
  assign after_write$060 = after_write[ 60];
  assign after_write$061 = after_write[ 61];
  assign after_write$062 = after_write[ 62];
  logic    [   0:0] regs[0:62];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  assign regs$002 = regs[  2];
  assign regs$003 = regs[  3];
  assign regs$004 = regs[  4];
  assign regs$005 = regs[  5];
  assign regs$006 = regs[  6];
  assign regs$007 = regs[  7];
  assign regs$008 = regs[  8];
  assign regs$009 = regs[  9];
  assign regs$010 = regs[ 10];
  assign regs$011 = regs[ 11];
  assign regs$012 = regs[ 12];
  assign regs$013 = regs[ 13];
  assign regs$014 = regs[ 14];
  assign regs$015 = regs[ 15];
  assign regs$016 = regs[ 16];
  assign regs$017 = regs[ 17];
  assign regs$018 = regs[ 18];
  assign regs$019 = regs[ 19];
  assign regs$020 = regs[ 20];
  assign regs$021 = regs[ 21];
  assign regs$022 = regs[ 22];
  assign regs$023 = regs[ 23];
  assign regs$024 = regs[ 24];
  assign regs$025 = regs[ 25];
  assign regs$026 = regs[ 26];
  assign regs$027 = regs[ 27];
  assign regs$028 = regs[ 28];
  assign regs$029 = regs[ 29];
  assign regs$030 = regs[ 30];
  assign regs$031 = regs[ 31];
  assign regs$032 = regs[ 32];
  assign regs$033 = regs[ 33];
  assign regs$034 = regs[ 34];
  assign regs$035 = regs[ 35];
  assign regs$036 = regs[ 36];
  assign regs$037 = regs[ 37];
  assign regs$038 = regs[ 38];
  assign regs$039 = regs[ 39];
  assign regs$040 = regs[ 40];
  assign regs$041 = regs[ 41];
  assign regs$042 = regs[ 42];
  assign regs$043 = regs[ 43];
  assign regs$044 = regs[ 44];
  assign regs$045 = regs[ 45];
  assign regs$046 = regs[ 46];
  assign regs$047 = regs[ 47];
  assign regs$048 = regs[ 48];
  assign regs$049 = regs[ 49];
  assign regs$050 = regs[ 50];
  assign regs$051 = regs[ 51];
  assign regs$052 = regs[ 52];
  assign regs$053 = regs[ 53];
  assign regs$054 = regs[ 54];
  assign regs$055 = regs[ 55];
  assign regs$056 = regs[ 56];
  assign regs$057 = regs[ 57];
  assign regs$058 = regs[ 58];
  assign regs$059 = regs[ 59];
  assign regs$060 = regs[ 60];
  assign regs$061 = regs[ 61];
  assign regs$062 = regs[ 62];
  logic   [   0:0] set_in_[0:62];
  assign set_in_[  0] = set_in_$000;
  assign set_in_[  1] = set_in_$001;
  assign set_in_[  2] = set_in_$002;
  assign set_in_[  3] = set_in_$003;
  assign set_in_[  4] = set_in_$004;
  assign set_in_[  5] = set_in_$005;
  assign set_in_[  6] = set_in_$006;
  assign set_in_[  7] = set_in_$007;
  assign set_in_[  8] = set_in_$008;
  assign set_in_[  9] = set_in_$009;
  assign set_in_[ 10] = set_in_$010;
  assign set_in_[ 11] = set_in_$011;
  assign set_in_[ 12] = set_in_$012;
  assign set_in_[ 13] = set_in_$013;
  assign set_in_[ 14] = set_in_$014;
  assign set_in_[ 15] = set_in_$015;
  assign set_in_[ 16] = set_in_$016;
  assign set_in_[ 17] = set_in_$017;
  assign set_in_[ 18] = set_in_$018;
  assign set_in_[ 19] = set_in_$019;
  assign set_in_[ 20] = set_in_$020;
  assign set_in_[ 21] = set_in_$021;
  assign set_in_[ 22] = set_in_$022;
  assign set_in_[ 23] = set_in_$023;
  assign set_in_[ 24] = set_in_$024;
  assign set_in_[ 25] = set_in_$025;
  assign set_in_[ 26] = set_in_$026;
  assign set_in_[ 27] = set_in_$027;
  assign set_in_[ 28] = set_in_$028;
  assign set_in_[ 29] = set_in_$029;
  assign set_in_[ 30] = set_in_$030;
  assign set_in_[ 31] = set_in_$031;
  assign set_in_[ 32] = set_in_$032;
  assign set_in_[ 33] = set_in_$033;
  assign set_in_[ 34] = set_in_$034;
  assign set_in_[ 35] = set_in_$035;
  assign set_in_[ 36] = set_in_$036;
  assign set_in_[ 37] = set_in_$037;
  assign set_in_[ 38] = set_in_$038;
  assign set_in_[ 39] = set_in_$039;
  assign set_in_[ 40] = set_in_$040;
  assign set_in_[ 41] = set_in_$041;
  assign set_in_[ 42] = set_in_$042;
  assign set_in_[ 43] = set_in_$043;
  assign set_in_[ 44] = set_in_$044;
  assign set_in_[ 45] = set_in_$045;
  assign set_in_[ 46] = set_in_$046;
  assign set_in_[ 47] = set_in_$047;
  assign set_in_[ 48] = set_in_$048;
  assign set_in_[ 49] = set_in_$049;
  assign set_in_[ 50] = set_in_$050;
  assign set_in_[ 51] = set_in_$051;
  assign set_in_[ 52] = set_in_$052;
  assign set_in_[ 53] = set_in_$053;
  assign set_in_[ 54] = set_in_$054;
  assign set_in_[ 55] = set_in_$055;
  assign set_in_[ 56] = set_in_$056;
  assign set_in_[ 57] = set_in_$057;
  assign set_in_[ 58] = set_in_$058;
  assign set_in_[ 59] = set_in_$059;
  assign set_in_[ 60] = set_in_$060;
  assign set_in_[ 61] = set_in_$061;
  assign set_in_[ 62] = set_in_$062;
  logic   [   5:0] write_addr[0:1];
  assign write_addr[  0] = write_addr$000;
  assign write_addr[  1] = write_addr$001;
  logic   [   0:0] write_call[0:1];
  assign write_call[  0] = write_call$000;
  assign write_call[  1] = write_call$001;
  logic   [   0:0] write_data[0:1];
  assign write_data[  0] = write_data$000;
  assign write_data[  1] = write_data$001;
  logic    [   0:0] write_inc[0:125];
  assign write_inc$000 = write_inc[  0];
  assign write_inc$001 = write_inc[  1];
  assign write_inc$002 = write_inc[  2];
  assign write_inc$003 = write_inc[  3];
  assign write_inc$004 = write_inc[  4];
  assign write_inc$005 = write_inc[  5];
  assign write_inc$006 = write_inc[  6];
  assign write_inc$007 = write_inc[  7];
  assign write_inc$008 = write_inc[  8];
  assign write_inc$009 = write_inc[  9];
  assign write_inc$010 = write_inc[ 10];
  assign write_inc$011 = write_inc[ 11];
  assign write_inc$012 = write_inc[ 12];
  assign write_inc$013 = write_inc[ 13];
  assign write_inc$014 = write_inc[ 14];
  assign write_inc$015 = write_inc[ 15];
  assign write_inc$016 = write_inc[ 16];
  assign write_inc$017 = write_inc[ 17];
  assign write_inc$018 = write_inc[ 18];
  assign write_inc$019 = write_inc[ 19];
  assign write_inc$020 = write_inc[ 20];
  assign write_inc$021 = write_inc[ 21];
  assign write_inc$022 = write_inc[ 22];
  assign write_inc$023 = write_inc[ 23];
  assign write_inc$024 = write_inc[ 24];
  assign write_inc$025 = write_inc[ 25];
  assign write_inc$026 = write_inc[ 26];
  assign write_inc$027 = write_inc[ 27];
  assign write_inc$028 = write_inc[ 28];
  assign write_inc$029 = write_inc[ 29];
  assign write_inc$030 = write_inc[ 30];
  assign write_inc$031 = write_inc[ 31];
  assign write_inc$032 = write_inc[ 32];
  assign write_inc$033 = write_inc[ 33];
  assign write_inc$034 = write_inc[ 34];
  assign write_inc$035 = write_inc[ 35];
  assign write_inc$036 = write_inc[ 36];
  assign write_inc$037 = write_inc[ 37];
  assign write_inc$038 = write_inc[ 38];
  assign write_inc$039 = write_inc[ 39];
  assign write_inc$040 = write_inc[ 40];
  assign write_inc$041 = write_inc[ 41];
  assign write_inc$042 = write_inc[ 42];
  assign write_inc$043 = write_inc[ 43];
  assign write_inc$044 = write_inc[ 44];
  assign write_inc$045 = write_inc[ 45];
  assign write_inc$046 = write_inc[ 46];
  assign write_inc$047 = write_inc[ 47];
  assign write_inc$048 = write_inc[ 48];
  assign write_inc$049 = write_inc[ 49];
  assign write_inc$050 = write_inc[ 50];
  assign write_inc$051 = write_inc[ 51];
  assign write_inc$052 = write_inc[ 52];
  assign write_inc$053 = write_inc[ 53];
  assign write_inc$054 = write_inc[ 54];
  assign write_inc$055 = write_inc[ 55];
  assign write_inc$056 = write_inc[ 56];
  assign write_inc$057 = write_inc[ 57];
  assign write_inc$058 = write_inc[ 58];
  assign write_inc$059 = write_inc[ 59];
  assign write_inc$060 = write_inc[ 60];
  assign write_inc$061 = write_inc[ 61];
  assign write_inc$062 = write_inc[ 62];
  assign write_inc$063 = write_inc[ 63];
  assign write_inc$064 = write_inc[ 64];
  assign write_inc$065 = write_inc[ 65];
  assign write_inc$066 = write_inc[ 66];
  assign write_inc$067 = write_inc[ 67];
  assign write_inc$068 = write_inc[ 68];
  assign write_inc$069 = write_inc[ 69];
  assign write_inc$070 = write_inc[ 70];
  assign write_inc$071 = write_inc[ 71];
  assign write_inc$072 = write_inc[ 72];
  assign write_inc$073 = write_inc[ 73];
  assign write_inc$074 = write_inc[ 74];
  assign write_inc$075 = write_inc[ 75];
  assign write_inc$076 = write_inc[ 76];
  assign write_inc$077 = write_inc[ 77];
  assign write_inc$078 = write_inc[ 78];
  assign write_inc$079 = write_inc[ 79];
  assign write_inc$080 = write_inc[ 80];
  assign write_inc$081 = write_inc[ 81];
  assign write_inc$082 = write_inc[ 82];
  assign write_inc$083 = write_inc[ 83];
  assign write_inc$084 = write_inc[ 84];
  assign write_inc$085 = write_inc[ 85];
  assign write_inc$086 = write_inc[ 86];
  assign write_inc$087 = write_inc[ 87];
  assign write_inc$088 = write_inc[ 88];
  assign write_inc$089 = write_inc[ 89];
  assign write_inc$090 = write_inc[ 90];
  assign write_inc$091 = write_inc[ 91];
  assign write_inc$092 = write_inc[ 92];
  assign write_inc$093 = write_inc[ 93];
  assign write_inc$094 = write_inc[ 94];
  assign write_inc$095 = write_inc[ 95];
  assign write_inc$096 = write_inc[ 96];
  assign write_inc$097 = write_inc[ 97];
  assign write_inc$098 = write_inc[ 98];
  assign write_inc$099 = write_inc[ 99];
  assign write_inc$100 = write_inc[100];
  assign write_inc$101 = write_inc[101];
  assign write_inc$102 = write_inc[102];
  assign write_inc$103 = write_inc[103];
  assign write_inc$104 = write_inc[104];
  assign write_inc$105 = write_inc[105];
  assign write_inc$106 = write_inc[106];
  assign write_inc$107 = write_inc[107];
  assign write_inc$108 = write_inc[108];
  assign write_inc$109 = write_inc[109];
  assign write_inc$110 = write_inc[110];
  assign write_inc$111 = write_inc[111];
  assign write_inc$112 = write_inc[112];
  assign write_inc$113 = write_inc[113];
  assign write_inc$114 = write_inc[114];
  assign write_inc$115 = write_inc[115];
  assign write_inc$116 = write_inc[116];
  assign write_inc$117 = write_inc[117];
  assign write_inc$118 = write_inc[118];
  assign write_inc$119 = write_inc[119];
  assign write_inc$120 = write_inc[120];
  assign write_inc$121 = write_inc[121];
  assign write_inc$122 = write_inc[122];
  assign write_inc$123 = write_inc[123];
  assign write_inc$124 = write_inc[124];
  assign write_inc$125 = write_inc[125];

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[0] <= 1;
    end
    else begin
      regs[0] <= after_set[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[1] <= 1;
    end
    else begin
      regs[1] <= after_set[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[2] <= 1;
    end
    else begin
      regs[2] <= after_set[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[3] <= 1;
    end
    else begin
      regs[3] <= after_set[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[4] <= 1;
    end
    else begin
      regs[4] <= after_set[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[5] <= 1;
    end
    else begin
      regs[5] <= after_set[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[6] <= 1;
    end
    else begin
      regs[6] <= after_set[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[7] <= 1;
    end
    else begin
      regs[7] <= after_set[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[8] <= 1;
    end
    else begin
      regs[8] <= after_set[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[9] <= 1;
    end
    else begin
      regs[9] <= after_set[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[10] <= 1;
    end
    else begin
      regs[10] <= after_set[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[11] <= 1;
    end
    else begin
      regs[11] <= after_set[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[12] <= 1;
    end
    else begin
      regs[12] <= after_set[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[13] <= 1;
    end
    else begin
      regs[13] <= after_set[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[14] <= 1;
    end
    else begin
      regs[14] <= after_set[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[15] <= 1;
    end
    else begin
      regs[15] <= after_set[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[16] <= 1;
    end
    else begin
      regs[16] <= after_set[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[17] <= 1;
    end
    else begin
      regs[17] <= after_set[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[18] <= 1;
    end
    else begin
      regs[18] <= after_set[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[19] <= 1;
    end
    else begin
      regs[19] <= after_set[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[20] <= 1;
    end
    else begin
      regs[20] <= after_set[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[21] <= 1;
    end
    else begin
      regs[21] <= after_set[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[22] <= 1;
    end
    else begin
      regs[22] <= after_set[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[23] <= 1;
    end
    else begin
      regs[23] <= after_set[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[24] <= 1;
    end
    else begin
      regs[24] <= after_set[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[25] <= 1;
    end
    else begin
      regs[25] <= after_set[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[26] <= 1;
    end
    else begin
      regs[26] <= after_set[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[27] <= 1;
    end
    else begin
      regs[27] <= after_set[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[28] <= 1;
    end
    else begin
      regs[28] <= after_set[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[29] <= 1;
    end
    else begin
      regs[29] <= after_set[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[30] <= 1;
    end
    else begin
      regs[30] <= after_set[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[31] <= 1;
    end
    else begin
      regs[31] <= after_set[31];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[32] <= 0;
    end
    else begin
      regs[32] <= after_set[32];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[33] <= 0;
    end
    else begin
      regs[33] <= after_set[33];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[34] <= 0;
    end
    else begin
      regs[34] <= after_set[34];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[35] <= 0;
    end
    else begin
      regs[35] <= after_set[35];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[36] <= 0;
    end
    else begin
      regs[36] <= after_set[36];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[37] <= 0;
    end
    else begin
      regs[37] <= after_set[37];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[38] <= 0;
    end
    else begin
      regs[38] <= after_set[38];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[39] <= 0;
    end
    else begin
      regs[39] <= after_set[39];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[40] <= 0;
    end
    else begin
      regs[40] <= after_set[40];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[41] <= 0;
    end
    else begin
      regs[41] <= after_set[41];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[42] <= 0;
    end
    else begin
      regs[42] <= after_set[42];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[43] <= 0;
    end
    else begin
      regs[43] <= after_set[43];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[44] <= 0;
    end
    else begin
      regs[44] <= after_set[44];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[45] <= 0;
    end
    else begin
      regs[45] <= after_set[45];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[46] <= 0;
    end
    else begin
      regs[46] <= after_set[46];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[47] <= 0;
    end
    else begin
      regs[47] <= after_set[47];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[48] <= 0;
    end
    else begin
      regs[48] <= after_set[48];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[49] <= 0;
    end
    else begin
      regs[49] <= after_set[49];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[50] <= 0;
    end
    else begin
      regs[50] <= after_set[50];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[51] <= 0;
    end
    else begin
      regs[51] <= after_set[51];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[52] <= 0;
    end
    else begin
      regs[52] <= after_set[52];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[53] <= 0;
    end
    else begin
      regs[53] <= after_set[53];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[54] <= 0;
    end
    else begin
      regs[54] <= after_set[54];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[55] <= 0;
    end
    else begin
      regs[55] <= after_set[55];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[56] <= 0;
    end
    else begin
      regs[56] <= after_set[56];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[57] <= 0;
    end
    else begin
      regs[57] <= after_set[57];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[58] <= 0;
    end
    else begin
      regs[58] <= after_set[58];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[59] <= 0;
    end
    else begin
      regs[59] <= after_set[59];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[60] <= 0;
    end
    else begin
      regs[60] <= after_set[60];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[61] <= 0;
    end
    else begin
      regs[61] <= after_set[61];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[62] <= 0;
    end
    else begin
      regs[62] <= after_set[62];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 0))) begin
      write_inc[0] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[0] = regs[0];
      end
      else begin
        write_inc[0] = write_inc[-63];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 0))) begin
      write_inc[63] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[63] = regs[0];
      end
      else begin
        write_inc[63] = write_inc[0];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[0] = write_inc[63];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[0] = set_in_[0];
    end
    else begin
      after_set[0] = after_write[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 1))) begin
      write_inc[1] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[1] = regs[1];
      end
      else begin
        write_inc[1] = write_inc[-62];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 1))) begin
      write_inc[64] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[64] = regs[1];
      end
      else begin
        write_inc[64] = write_inc[1];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[1] = write_inc[64];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[1] = set_in_[1];
    end
    else begin
      after_set[1] = after_write[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 2))) begin
      write_inc[2] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[2] = regs[2];
      end
      else begin
        write_inc[2] = write_inc[-61];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 2))) begin
      write_inc[65] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[65] = regs[2];
      end
      else begin
        write_inc[65] = write_inc[2];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[2] = write_inc[65];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[2] = set_in_[2];
    end
    else begin
      after_set[2] = after_write[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 3))) begin
      write_inc[3] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[3] = regs[3];
      end
      else begin
        write_inc[3] = write_inc[-60];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 3))) begin
      write_inc[66] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[66] = regs[3];
      end
      else begin
        write_inc[66] = write_inc[3];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[3] = write_inc[66];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[3] = set_in_[3];
    end
    else begin
      after_set[3] = after_write[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 4))) begin
      write_inc[4] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[4] = regs[4];
      end
      else begin
        write_inc[4] = write_inc[-59];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 4))) begin
      write_inc[67] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[67] = regs[4];
      end
      else begin
        write_inc[67] = write_inc[4];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[4] = write_inc[67];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[4] = set_in_[4];
    end
    else begin
      after_set[4] = after_write[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 5))) begin
      write_inc[5] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[5] = regs[5];
      end
      else begin
        write_inc[5] = write_inc[-58];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 5))) begin
      write_inc[68] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[68] = regs[5];
      end
      else begin
        write_inc[68] = write_inc[5];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[5] = write_inc[68];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[5] = set_in_[5];
    end
    else begin
      after_set[5] = after_write[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 6))) begin
      write_inc[6] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[6] = regs[6];
      end
      else begin
        write_inc[6] = write_inc[-57];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 6))) begin
      write_inc[69] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[69] = regs[6];
      end
      else begin
        write_inc[69] = write_inc[6];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[6] = write_inc[69];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[6] = set_in_[6];
    end
    else begin
      after_set[6] = after_write[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 7))) begin
      write_inc[7] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[7] = regs[7];
      end
      else begin
        write_inc[7] = write_inc[-56];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 7))) begin
      write_inc[70] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[70] = regs[7];
      end
      else begin
        write_inc[70] = write_inc[7];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[7] = write_inc[70];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[7] = set_in_[7];
    end
    else begin
      after_set[7] = after_write[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 8))) begin
      write_inc[8] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[8] = regs[8];
      end
      else begin
        write_inc[8] = write_inc[-55];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 8))) begin
      write_inc[71] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[71] = regs[8];
      end
      else begin
        write_inc[71] = write_inc[8];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[8] = write_inc[71];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[8] = set_in_[8];
    end
    else begin
      after_set[8] = after_write[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 9))) begin
      write_inc[9] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[9] = regs[9];
      end
      else begin
        write_inc[9] = write_inc[-54];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 9))) begin
      write_inc[72] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[72] = regs[9];
      end
      else begin
        write_inc[72] = write_inc[9];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[9] = write_inc[72];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[9] = set_in_[9];
    end
    else begin
      after_set[9] = after_write[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 10))) begin
      write_inc[10] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[10] = regs[10];
      end
      else begin
        write_inc[10] = write_inc[-53];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 10))) begin
      write_inc[73] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[73] = regs[10];
      end
      else begin
        write_inc[73] = write_inc[10];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[10] = write_inc[73];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[10] = set_in_[10];
    end
    else begin
      after_set[10] = after_write[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 11))) begin
      write_inc[11] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[11] = regs[11];
      end
      else begin
        write_inc[11] = write_inc[-52];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 11))) begin
      write_inc[74] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[74] = regs[11];
      end
      else begin
        write_inc[74] = write_inc[11];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[11] = write_inc[74];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[11] = set_in_[11];
    end
    else begin
      after_set[11] = after_write[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 12))) begin
      write_inc[12] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[12] = regs[12];
      end
      else begin
        write_inc[12] = write_inc[-51];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 12))) begin
      write_inc[75] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[75] = regs[12];
      end
      else begin
        write_inc[75] = write_inc[12];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[12] = write_inc[75];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[12] = set_in_[12];
    end
    else begin
      after_set[12] = after_write[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 13))) begin
      write_inc[13] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[13] = regs[13];
      end
      else begin
        write_inc[13] = write_inc[-50];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 13))) begin
      write_inc[76] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[76] = regs[13];
      end
      else begin
        write_inc[76] = write_inc[13];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[13] = write_inc[76];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[13] = set_in_[13];
    end
    else begin
      after_set[13] = after_write[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 14))) begin
      write_inc[14] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[14] = regs[14];
      end
      else begin
        write_inc[14] = write_inc[-49];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 14))) begin
      write_inc[77] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[77] = regs[14];
      end
      else begin
        write_inc[77] = write_inc[14];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[14] = write_inc[77];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[14] = set_in_[14];
    end
    else begin
      after_set[14] = after_write[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 15))) begin
      write_inc[15] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[15] = regs[15];
      end
      else begin
        write_inc[15] = write_inc[-48];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 15))) begin
      write_inc[78] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[78] = regs[15];
      end
      else begin
        write_inc[78] = write_inc[15];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[15] = write_inc[78];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[15] = set_in_[15];
    end
    else begin
      after_set[15] = after_write[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 16))) begin
      write_inc[16] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[16] = regs[16];
      end
      else begin
        write_inc[16] = write_inc[-47];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 16))) begin
      write_inc[79] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[79] = regs[16];
      end
      else begin
        write_inc[79] = write_inc[16];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[16] = write_inc[79];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[16] = set_in_[16];
    end
    else begin
      after_set[16] = after_write[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 17))) begin
      write_inc[17] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[17] = regs[17];
      end
      else begin
        write_inc[17] = write_inc[-46];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 17))) begin
      write_inc[80] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[80] = regs[17];
      end
      else begin
        write_inc[80] = write_inc[17];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[17] = write_inc[80];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[17] = set_in_[17];
    end
    else begin
      after_set[17] = after_write[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 18))) begin
      write_inc[18] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[18] = regs[18];
      end
      else begin
        write_inc[18] = write_inc[-45];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 18))) begin
      write_inc[81] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[81] = regs[18];
      end
      else begin
        write_inc[81] = write_inc[18];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[18] = write_inc[81];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[18] = set_in_[18];
    end
    else begin
      after_set[18] = after_write[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 19))) begin
      write_inc[19] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[19] = regs[19];
      end
      else begin
        write_inc[19] = write_inc[-44];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 19))) begin
      write_inc[82] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[82] = regs[19];
      end
      else begin
        write_inc[82] = write_inc[19];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[19] = write_inc[82];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[19] = set_in_[19];
    end
    else begin
      after_set[19] = after_write[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 20))) begin
      write_inc[20] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[20] = regs[20];
      end
      else begin
        write_inc[20] = write_inc[-43];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 20))) begin
      write_inc[83] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[83] = regs[20];
      end
      else begin
        write_inc[83] = write_inc[20];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[20] = write_inc[83];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[20] = set_in_[20];
    end
    else begin
      after_set[20] = after_write[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 21))) begin
      write_inc[21] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[21] = regs[21];
      end
      else begin
        write_inc[21] = write_inc[-42];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 21))) begin
      write_inc[84] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[84] = regs[21];
      end
      else begin
        write_inc[84] = write_inc[21];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[21] = write_inc[84];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[21] = set_in_[21];
    end
    else begin
      after_set[21] = after_write[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 22))) begin
      write_inc[22] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[22] = regs[22];
      end
      else begin
        write_inc[22] = write_inc[-41];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 22))) begin
      write_inc[85] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[85] = regs[22];
      end
      else begin
        write_inc[85] = write_inc[22];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[22] = write_inc[85];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[22] = set_in_[22];
    end
    else begin
      after_set[22] = after_write[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 23))) begin
      write_inc[23] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[23] = regs[23];
      end
      else begin
        write_inc[23] = write_inc[-40];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 23))) begin
      write_inc[86] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[86] = regs[23];
      end
      else begin
        write_inc[86] = write_inc[23];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[23] = write_inc[86];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[23] = set_in_[23];
    end
    else begin
      after_set[23] = after_write[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 24))) begin
      write_inc[24] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[24] = regs[24];
      end
      else begin
        write_inc[24] = write_inc[-39];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 24))) begin
      write_inc[87] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[87] = regs[24];
      end
      else begin
        write_inc[87] = write_inc[24];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[24] = write_inc[87];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[24] = set_in_[24];
    end
    else begin
      after_set[24] = after_write[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 25))) begin
      write_inc[25] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[25] = regs[25];
      end
      else begin
        write_inc[25] = write_inc[-38];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 25))) begin
      write_inc[88] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[88] = regs[25];
      end
      else begin
        write_inc[88] = write_inc[25];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[25] = write_inc[88];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[25] = set_in_[25];
    end
    else begin
      after_set[25] = after_write[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 26))) begin
      write_inc[26] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[26] = regs[26];
      end
      else begin
        write_inc[26] = write_inc[-37];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 26))) begin
      write_inc[89] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[89] = regs[26];
      end
      else begin
        write_inc[89] = write_inc[26];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[26] = write_inc[89];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[26] = set_in_[26];
    end
    else begin
      after_set[26] = after_write[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 27))) begin
      write_inc[27] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[27] = regs[27];
      end
      else begin
        write_inc[27] = write_inc[-36];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 27))) begin
      write_inc[90] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[90] = regs[27];
      end
      else begin
        write_inc[90] = write_inc[27];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[27] = write_inc[90];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[27] = set_in_[27];
    end
    else begin
      after_set[27] = after_write[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 28))) begin
      write_inc[28] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[28] = regs[28];
      end
      else begin
        write_inc[28] = write_inc[-35];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 28))) begin
      write_inc[91] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[91] = regs[28];
      end
      else begin
        write_inc[91] = write_inc[28];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[28] = write_inc[91];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[28] = set_in_[28];
    end
    else begin
      after_set[28] = after_write[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 29))) begin
      write_inc[29] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[29] = regs[29];
      end
      else begin
        write_inc[29] = write_inc[-34];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 29))) begin
      write_inc[92] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[92] = regs[29];
      end
      else begin
        write_inc[92] = write_inc[29];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[29] = write_inc[92];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[29] = set_in_[29];
    end
    else begin
      after_set[29] = after_write[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 30))) begin
      write_inc[30] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[30] = regs[30];
      end
      else begin
        write_inc[30] = write_inc[-33];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 30))) begin
      write_inc[93] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[93] = regs[30];
      end
      else begin
        write_inc[93] = write_inc[30];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[30] = write_inc[93];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[30] = set_in_[30];
    end
    else begin
      after_set[30] = after_write[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 31))) begin
      write_inc[31] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[31] = regs[31];
      end
      else begin
        write_inc[31] = write_inc[-32];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 31))) begin
      write_inc[94] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[94] = regs[31];
      end
      else begin
        write_inc[94] = write_inc[31];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[31] = write_inc[94];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[31] = set_in_[31];
    end
    else begin
      after_set[31] = after_write[31];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 32))) begin
      write_inc[32] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[32] = regs[32];
      end
      else begin
        write_inc[32] = write_inc[-31];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 32))) begin
      write_inc[95] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[95] = regs[32];
      end
      else begin
        write_inc[95] = write_inc[32];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[32] = write_inc[95];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[32] = set_in_[32];
    end
    else begin
      after_set[32] = after_write[32];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 33))) begin
      write_inc[33] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[33] = regs[33];
      end
      else begin
        write_inc[33] = write_inc[-30];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 33))) begin
      write_inc[96] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[96] = regs[33];
      end
      else begin
        write_inc[96] = write_inc[33];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[33] = write_inc[96];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[33] = set_in_[33];
    end
    else begin
      after_set[33] = after_write[33];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 34))) begin
      write_inc[34] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[34] = regs[34];
      end
      else begin
        write_inc[34] = write_inc[-29];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 34))) begin
      write_inc[97] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[97] = regs[34];
      end
      else begin
        write_inc[97] = write_inc[34];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[34] = write_inc[97];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[34] = set_in_[34];
    end
    else begin
      after_set[34] = after_write[34];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 35))) begin
      write_inc[35] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[35] = regs[35];
      end
      else begin
        write_inc[35] = write_inc[-28];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 35))) begin
      write_inc[98] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[98] = regs[35];
      end
      else begin
        write_inc[98] = write_inc[35];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[35] = write_inc[98];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[35] = set_in_[35];
    end
    else begin
      after_set[35] = after_write[35];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 36))) begin
      write_inc[36] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[36] = regs[36];
      end
      else begin
        write_inc[36] = write_inc[-27];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 36))) begin
      write_inc[99] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[99] = regs[36];
      end
      else begin
        write_inc[99] = write_inc[36];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[36] = write_inc[99];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[36] = set_in_[36];
    end
    else begin
      after_set[36] = after_write[36];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 37))) begin
      write_inc[37] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[37] = regs[37];
      end
      else begin
        write_inc[37] = write_inc[-26];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 37))) begin
      write_inc[100] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[100] = regs[37];
      end
      else begin
        write_inc[100] = write_inc[37];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[37] = write_inc[100];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[37] = set_in_[37];
    end
    else begin
      after_set[37] = after_write[37];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 38))) begin
      write_inc[38] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[38] = regs[38];
      end
      else begin
        write_inc[38] = write_inc[-25];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 38))) begin
      write_inc[101] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[101] = regs[38];
      end
      else begin
        write_inc[101] = write_inc[38];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[38] = write_inc[101];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[38] = set_in_[38];
    end
    else begin
      after_set[38] = after_write[38];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 39))) begin
      write_inc[39] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[39] = regs[39];
      end
      else begin
        write_inc[39] = write_inc[-24];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 39))) begin
      write_inc[102] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[102] = regs[39];
      end
      else begin
        write_inc[102] = write_inc[39];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[39] = write_inc[102];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[39] = set_in_[39];
    end
    else begin
      after_set[39] = after_write[39];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 40))) begin
      write_inc[40] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[40] = regs[40];
      end
      else begin
        write_inc[40] = write_inc[-23];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 40))) begin
      write_inc[103] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[103] = regs[40];
      end
      else begin
        write_inc[103] = write_inc[40];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[40] = write_inc[103];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[40] = set_in_[40];
    end
    else begin
      after_set[40] = after_write[40];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 41))) begin
      write_inc[41] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[41] = regs[41];
      end
      else begin
        write_inc[41] = write_inc[-22];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 41))) begin
      write_inc[104] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[104] = regs[41];
      end
      else begin
        write_inc[104] = write_inc[41];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[41] = write_inc[104];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[41] = set_in_[41];
    end
    else begin
      after_set[41] = after_write[41];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 42))) begin
      write_inc[42] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[42] = regs[42];
      end
      else begin
        write_inc[42] = write_inc[-21];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 42))) begin
      write_inc[105] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[105] = regs[42];
      end
      else begin
        write_inc[105] = write_inc[42];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[42] = write_inc[105];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[42] = set_in_[42];
    end
    else begin
      after_set[42] = after_write[42];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 43))) begin
      write_inc[43] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[43] = regs[43];
      end
      else begin
        write_inc[43] = write_inc[-20];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 43))) begin
      write_inc[106] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[106] = regs[43];
      end
      else begin
        write_inc[106] = write_inc[43];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[43] = write_inc[106];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[43] = set_in_[43];
    end
    else begin
      after_set[43] = after_write[43];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 44))) begin
      write_inc[44] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[44] = regs[44];
      end
      else begin
        write_inc[44] = write_inc[-19];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 44))) begin
      write_inc[107] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[107] = regs[44];
      end
      else begin
        write_inc[107] = write_inc[44];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[44] = write_inc[107];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[44] = set_in_[44];
    end
    else begin
      after_set[44] = after_write[44];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 45))) begin
      write_inc[45] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[45] = regs[45];
      end
      else begin
        write_inc[45] = write_inc[-18];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 45))) begin
      write_inc[108] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[108] = regs[45];
      end
      else begin
        write_inc[108] = write_inc[45];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[45] = write_inc[108];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[45] = set_in_[45];
    end
    else begin
      after_set[45] = after_write[45];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 46))) begin
      write_inc[46] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[46] = regs[46];
      end
      else begin
        write_inc[46] = write_inc[-17];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 46))) begin
      write_inc[109] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[109] = regs[46];
      end
      else begin
        write_inc[109] = write_inc[46];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[46] = write_inc[109];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[46] = set_in_[46];
    end
    else begin
      after_set[46] = after_write[46];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 47))) begin
      write_inc[47] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[47] = regs[47];
      end
      else begin
        write_inc[47] = write_inc[-16];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 47))) begin
      write_inc[110] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[110] = regs[47];
      end
      else begin
        write_inc[110] = write_inc[47];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[47] = write_inc[110];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[47] = set_in_[47];
    end
    else begin
      after_set[47] = after_write[47];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 48))) begin
      write_inc[48] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[48] = regs[48];
      end
      else begin
        write_inc[48] = write_inc[-15];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 48))) begin
      write_inc[111] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[111] = regs[48];
      end
      else begin
        write_inc[111] = write_inc[48];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[48] = write_inc[111];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[48] = set_in_[48];
    end
    else begin
      after_set[48] = after_write[48];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 49))) begin
      write_inc[49] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[49] = regs[49];
      end
      else begin
        write_inc[49] = write_inc[-14];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 49))) begin
      write_inc[112] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[112] = regs[49];
      end
      else begin
        write_inc[112] = write_inc[49];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[49] = write_inc[112];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[49] = set_in_[49];
    end
    else begin
      after_set[49] = after_write[49];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 50))) begin
      write_inc[50] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[50] = regs[50];
      end
      else begin
        write_inc[50] = write_inc[-13];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 50))) begin
      write_inc[113] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[113] = regs[50];
      end
      else begin
        write_inc[113] = write_inc[50];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[50] = write_inc[113];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[50] = set_in_[50];
    end
    else begin
      after_set[50] = after_write[50];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 51))) begin
      write_inc[51] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[51] = regs[51];
      end
      else begin
        write_inc[51] = write_inc[-12];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 51))) begin
      write_inc[114] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[114] = regs[51];
      end
      else begin
        write_inc[114] = write_inc[51];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[51] = write_inc[114];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[51] = set_in_[51];
    end
    else begin
      after_set[51] = after_write[51];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 52))) begin
      write_inc[52] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[52] = regs[52];
      end
      else begin
        write_inc[52] = write_inc[-11];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 52))) begin
      write_inc[115] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[115] = regs[52];
      end
      else begin
        write_inc[115] = write_inc[52];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[52] = write_inc[115];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[52] = set_in_[52];
    end
    else begin
      after_set[52] = after_write[52];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 53))) begin
      write_inc[53] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[53] = regs[53];
      end
      else begin
        write_inc[53] = write_inc[-10];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 53))) begin
      write_inc[116] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[116] = regs[53];
      end
      else begin
        write_inc[116] = write_inc[53];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[53] = write_inc[116];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[53] = set_in_[53];
    end
    else begin
      after_set[53] = after_write[53];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 54))) begin
      write_inc[54] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[54] = regs[54];
      end
      else begin
        write_inc[54] = write_inc[-9];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 54))) begin
      write_inc[117] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[117] = regs[54];
      end
      else begin
        write_inc[117] = write_inc[54];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[54] = write_inc[117];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[54] = set_in_[54];
    end
    else begin
      after_set[54] = after_write[54];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 55))) begin
      write_inc[55] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[55] = regs[55];
      end
      else begin
        write_inc[55] = write_inc[-8];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 55))) begin
      write_inc[118] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[118] = regs[55];
      end
      else begin
        write_inc[118] = write_inc[55];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[55] = write_inc[118];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[55] = set_in_[55];
    end
    else begin
      after_set[55] = after_write[55];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 56))) begin
      write_inc[56] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[56] = regs[56];
      end
      else begin
        write_inc[56] = write_inc[-7];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 56))) begin
      write_inc[119] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[119] = regs[56];
      end
      else begin
        write_inc[119] = write_inc[56];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[56] = write_inc[119];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[56] = set_in_[56];
    end
    else begin
      after_set[56] = after_write[56];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 57))) begin
      write_inc[57] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[57] = regs[57];
      end
      else begin
        write_inc[57] = write_inc[-6];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 57))) begin
      write_inc[120] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[120] = regs[57];
      end
      else begin
        write_inc[120] = write_inc[57];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[57] = write_inc[120];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[57] = set_in_[57];
    end
    else begin
      after_set[57] = after_write[57];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 58))) begin
      write_inc[58] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[58] = regs[58];
      end
      else begin
        write_inc[58] = write_inc[-5];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 58))) begin
      write_inc[121] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[121] = regs[58];
      end
      else begin
        write_inc[121] = write_inc[58];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[58] = write_inc[121];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[58] = set_in_[58];
    end
    else begin
      after_set[58] = after_write[58];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 59))) begin
      write_inc[59] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[59] = regs[59];
      end
      else begin
        write_inc[59] = write_inc[-4];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 59))) begin
      write_inc[122] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[122] = regs[59];
      end
      else begin
        write_inc[122] = write_inc[59];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[59] = write_inc[122];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[59] = set_in_[59];
    end
    else begin
      after_set[59] = after_write[59];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 60))) begin
      write_inc[60] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[60] = regs[60];
      end
      else begin
        write_inc[60] = write_inc[-3];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 60))) begin
      write_inc[123] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[123] = regs[60];
      end
      else begin
        write_inc[123] = write_inc[60];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[60] = write_inc[123];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[60] = set_in_[60];
    end
    else begin
      after_set[60] = after_write[60];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 61))) begin
      write_inc[61] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[61] = regs[61];
      end
      else begin
        write_inc[61] = write_inc[-2];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 61))) begin
      write_inc[124] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[124] = regs[61];
      end
      else begin
        write_inc[124] = write_inc[61];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[61] = write_inc[124];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[61] = set_in_[61];
    end
    else begin
      after_set[61] = after_write[61];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 62))) begin
      write_inc[62] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[62] = regs[62];
      end
      else begin
        write_inc[62] = write_inc[-1];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[1]&&(write_addr[1] == 62))) begin
      write_inc[125] = write_data[1];
    end
    else begin
      if ((1 == 0)) begin
        write_inc[125] = regs[62];
      end
      else begin
        write_inc[125] = write_inc[62];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[62] = write_inc[125];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[62] = set_in_[62];
    end
    else begin
      after_set[62] = after_write[62];
    end
  end


endmodule // RegisterFile_0x39d647b3aea936a6

//-----------------------------------------------------------------------------
// Mux_0x1d47079284a028c3
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.mux {"dtype": 64, "nports": 2}
// PyMTL: verilator_xinit = zeros
module Mux_0x1d47079284a028c3
(
  input  logic [   0:0] clk,
  input  logic [  63:0] mux_in_$000,
  input  logic [  63:0] mux_in_$001,
  output logic  [  63:0] mux_out,
  input  logic [   0:0] mux_select,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nports = 2;


  // array declarations
  logic   [  63:0] mux_in_[0:1];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def select():
  //       assert s.mux_select < nports
  //       s.mux_out.v = s.mux_in_[s.mux_select]

  // logic for select()
  always @ (*) begin
    mux_out = mux_in_[mux_select];
  end


endmodule // Mux_0x1d47079284a028c3

//-----------------------------------------------------------------------------
// AsynchronousRAM_0xb915281a52f5e7
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.async_ram {"interface": "write[2] <C> (data: Bits(64), addr: Bits(6)) -> (); read[2] (addr: Bits(6)) -> (data: Bits(64))", "reset_values": 0}
// PyMTL: verilator_xinit = zeros
module AsynchronousRAM_0xb915281a52f5e7
(
  input  logic [   0:0] clk,
  input  logic [   5:0] read_addr$000,
  input  logic [   5:0] read_addr$001,
  output logic [  63:0] read_data$000,
  output logic [  63:0] read_data$001,
  input  logic [   0:0] reset,
  input  logic [   5:0] write_addr$000,
  input  logic [   5:0] write_addr$001,
  input  logic [   0:0] write_call$000,
  input  logic [   0:0] write_call$001,
  input  logic [  63:0] write_data$000,
  input  logic [  63:0] write_data$001
);

  // logic declarations
  logic   [  63:0] regs$000;
  logic   [  63:0] regs$001;
  logic   [  63:0] regs$002;
  logic   [  63:0] regs$003;
  logic   [  63:0] regs$004;
  logic   [  63:0] regs$005;
  logic   [  63:0] regs$006;
  logic   [  63:0] regs$007;
  logic   [  63:0] regs$008;
  logic   [  63:0] regs$009;
  logic   [  63:0] regs$010;
  logic   [  63:0] regs$011;
  logic   [  63:0] regs$012;
  logic   [  63:0] regs$013;
  logic   [  63:0] regs$014;
  logic   [  63:0] regs$015;
  logic   [  63:0] regs$016;
  logic   [  63:0] regs$017;
  logic   [  63:0] regs$018;
  logic   [  63:0] regs$019;
  logic   [  63:0] regs$020;
  logic   [  63:0] regs$021;
  logic   [  63:0] regs$022;
  logic   [  63:0] regs$023;
  logic   [  63:0] regs$024;
  logic   [  63:0] regs$025;
  logic   [  63:0] regs$026;
  logic   [  63:0] regs$027;
  logic   [  63:0] regs$028;
  logic   [  63:0] regs$029;
  logic   [  63:0] regs$030;
  logic   [  63:0] regs$031;
  logic   [  63:0] regs$032;
  logic   [  63:0] regs$033;
  logic   [  63:0] regs$034;
  logic   [  63:0] regs$035;
  logic   [  63:0] regs$036;
  logic   [  63:0] regs$037;
  logic   [  63:0] regs$038;
  logic   [  63:0] regs$039;
  logic   [  63:0] regs$040;
  logic   [  63:0] regs$041;
  logic   [  63:0] regs$042;
  logic   [  63:0] regs$043;
  logic   [  63:0] regs$044;
  logic   [  63:0] regs$045;
  logic   [  63:0] regs$046;
  logic   [  63:0] regs$047;
  logic   [  63:0] regs$048;
  logic   [  63:0] regs$049;
  logic   [  63:0] regs$050;
  logic   [  63:0] regs$051;
  logic   [  63:0] regs$052;
  logic   [  63:0] regs$053;
  logic   [  63:0] regs$054;
  logic   [  63:0] regs$055;
  logic   [  63:0] regs$056;
  logic   [  63:0] regs$057;
  logic   [  63:0] regs$058;
  logic   [  63:0] regs$059;
  logic   [  63:0] regs$060;
  logic   [  63:0] regs$061;
  logic   [  63:0] regs$062;
  logic   [  63:0] regs$063;


  // localparam declarations
  localparam num_read_ports = 2;
  localparam num_write_ports = 2;
  localparam nwords = 64;
  localparam reset_values = 0;

  // loop variable declarations
  integer i;
  integer j;


  // array declarations
  logic   [   5:0] read_addr[0:1];
  assign read_addr[  0] = read_addr$000;
  assign read_addr[  1] = read_addr$001;
  logic    [  63:0] read_data[0:1];
  assign read_data$000 = read_data[  0];
  assign read_data$001 = read_data[  1];
  logic    [  63:0] regs[0:63];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  assign regs$002 = regs[  2];
  assign regs$003 = regs[  3];
  assign regs$004 = regs[  4];
  assign regs$005 = regs[  5];
  assign regs$006 = regs[  6];
  assign regs$007 = regs[  7];
  assign regs$008 = regs[  8];
  assign regs$009 = regs[  9];
  assign regs$010 = regs[ 10];
  assign regs$011 = regs[ 11];
  assign regs$012 = regs[ 12];
  assign regs$013 = regs[ 13];
  assign regs$014 = regs[ 14];
  assign regs$015 = regs[ 15];
  assign regs$016 = regs[ 16];
  assign regs$017 = regs[ 17];
  assign regs$018 = regs[ 18];
  assign regs$019 = regs[ 19];
  assign regs$020 = regs[ 20];
  assign regs$021 = regs[ 21];
  assign regs$022 = regs[ 22];
  assign regs$023 = regs[ 23];
  assign regs$024 = regs[ 24];
  assign regs$025 = regs[ 25];
  assign regs$026 = regs[ 26];
  assign regs$027 = regs[ 27];
  assign regs$028 = regs[ 28];
  assign regs$029 = regs[ 29];
  assign regs$030 = regs[ 30];
  assign regs$031 = regs[ 31];
  assign regs$032 = regs[ 32];
  assign regs$033 = regs[ 33];
  assign regs$034 = regs[ 34];
  assign regs$035 = regs[ 35];
  assign regs$036 = regs[ 36];
  assign regs$037 = regs[ 37];
  assign regs$038 = regs[ 38];
  assign regs$039 = regs[ 39];
  assign regs$040 = regs[ 40];
  assign regs$041 = regs[ 41];
  assign regs$042 = regs[ 42];
  assign regs$043 = regs[ 43];
  assign regs$044 = regs[ 44];
  assign regs$045 = regs[ 45];
  assign regs$046 = regs[ 46];
  assign regs$047 = regs[ 47];
  assign regs$048 = regs[ 48];
  assign regs$049 = regs[ 49];
  assign regs$050 = regs[ 50];
  assign regs$051 = regs[ 51];
  assign regs$052 = regs[ 52];
  assign regs$053 = regs[ 53];
  assign regs$054 = regs[ 54];
  assign regs$055 = regs[ 55];
  assign regs$056 = regs[ 56];
  assign regs$057 = regs[ 57];
  assign regs$058 = regs[ 58];
  assign regs$059 = regs[ 59];
  assign regs$060 = regs[ 60];
  assign regs$061 = regs[ 61];
  assign regs$062 = regs[ 62];
  assign regs$063 = regs[ 63];
  logic   [   5:0] write_addr[0:1];
  assign write_addr[  0] = write_addr$000;
  assign write_addr[  1] = write_addr$001;
  logic   [   0:0] write_call[0:1];
  assign write_call[  0] = write_call$000;
  assign write_call[  1] = write_call$001;
  logic   [  63:0] write_data[0:1];
  assign write_data[  0] = write_data$000;
  assign write_data[  1] = write_data$001;

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def handle_writes():
  //         if s.reset:
  //           for i in range(nwords):
  //             s.regs[i].n = reset_values
  //         else:
  //           for i in range(num_write_ports):
  //             if s.write_call[i]:
  //               s.regs[s.write_addr[i]].n = s.write_data[i]

  // logic for handle_writes()
  always @ (posedge clk) begin
    if (reset) begin
      for (i=0; i < nwords; i=i+1)
      begin
        regs[i] <= reset_values;
      end
    end
    else begin
      for (i=0; i < num_write_ports; i=i+1)
      begin
        if (write_call[i]) begin
          regs[write_addr[i]] <= write_data[i];
        end
        else begin
        end
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_reads():
  //         for i in range(num_read_ports):
  //           s.read_data[i].v = s.regs[s.read_addr[i]]
  //           # Bypass logic
  //           for j in range(num_write_ports):
  //             if s.write_call[j] and s.write_addr[j] == s.read_addr[i]:
  //               s.read_data[i].v = s.write_data[j]

  // logic for handle_reads()
  always @ (*) begin
    for (i=0; i < num_read_ports; i=i+1)
    begin
      read_data[i] = regs[read_addr[i]];
      for (j=0; j < num_write_ports; j=j+1)
      begin
        if ((write_call[j]&&(write_addr[j] == read_addr[i]))) begin
          read_data[i] = write_data[j];
        end
        else begin
        end
      end
    end
  end


endmodule // AsynchronousRAM_0xb915281a52f5e7

//-----------------------------------------------------------------------------
// SnapshottingFreeList_0x68f914e32e2c4f6d
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.snapshotting_freelist {"freelist_impl": "<class 'util.rtl.freelist.FreeList'>", "nslots": 63, "nsnapshots": 2, "num_alloc_ports": 1, "num_free_ports": 2, "used_slots_initial": 31}
// PyMTL: verilator_xinit = zeros
module SnapshottingFreeList_0x68f914e32e2c4f6d
(
  input  logic [   0:0] alloc_call$000,
  output logic [   5:0] alloc_index$000,
  output logic [  62:0] alloc_mask$000,
  output logic [   0:0] alloc_rdy$000,
  input  logic [   0:0] clk,
  input  logic [   0:0] free_call$000,
  input  logic [   0:0] free_call$001,
  input  logic [   5:0] free_index$000,
  input  logic [   5:0] free_index$001,
  input  logic [   0:0] reset,
  input  logic [   0:0] reset_alloc_tracking_call,
  input  logic [   0:0] reset_alloc_tracking_target_id,
  input  logic [   0:0] revert_allocs_call,
  input  logic [   0:0] revert_allocs_source_id,
  input  logic [   0:0] set_call,
  input  logic [  62:0] set_state
);

  // register declarations
  logic    [   0:0] free_list$release_call;

  // snapshots$000 temporaries
  logic   [   0:0] snapshots$000$set_in_$000;
  logic   [   0:0] snapshots$000$set_in_$001;
  logic   [   0:0] snapshots$000$set_in_$002;
  logic   [   0:0] snapshots$000$set_in_$003;
  logic   [   0:0] snapshots$000$set_in_$004;
  logic   [   0:0] snapshots$000$set_in_$005;
  logic   [   0:0] snapshots$000$set_in_$006;
  logic   [   0:0] snapshots$000$set_in_$007;
  logic   [   0:0] snapshots$000$set_in_$008;
  logic   [   0:0] snapshots$000$set_in_$009;
  logic   [   0:0] snapshots$000$set_in_$010;
  logic   [   0:0] snapshots$000$set_in_$011;
  logic   [   0:0] snapshots$000$set_in_$012;
  logic   [   0:0] snapshots$000$set_in_$013;
  logic   [   0:0] snapshots$000$set_in_$014;
  logic   [   0:0] snapshots$000$set_in_$015;
  logic   [   0:0] snapshots$000$set_in_$016;
  logic   [   0:0] snapshots$000$set_in_$017;
  logic   [   0:0] snapshots$000$set_in_$018;
  logic   [   0:0] snapshots$000$set_in_$019;
  logic   [   0:0] snapshots$000$set_in_$020;
  logic   [   0:0] snapshots$000$set_in_$021;
  logic   [   0:0] snapshots$000$set_in_$022;
  logic   [   0:0] snapshots$000$set_in_$023;
  logic   [   0:0] snapshots$000$set_in_$024;
  logic   [   0:0] snapshots$000$set_in_$025;
  logic   [   0:0] snapshots$000$set_in_$026;
  logic   [   0:0] snapshots$000$set_in_$027;
  logic   [   0:0] snapshots$000$set_in_$028;
  logic   [   0:0] snapshots$000$set_in_$029;
  logic   [   0:0] snapshots$000$set_in_$030;
  logic   [   0:0] snapshots$000$set_in_$031;
  logic   [   0:0] snapshots$000$set_in_$032;
  logic   [   0:0] snapshots$000$set_in_$033;
  logic   [   0:0] snapshots$000$set_in_$034;
  logic   [   0:0] snapshots$000$set_in_$035;
  logic   [   0:0] snapshots$000$set_in_$036;
  logic   [   0:0] snapshots$000$set_in_$037;
  logic   [   0:0] snapshots$000$set_in_$038;
  logic   [   0:0] snapshots$000$set_in_$039;
  logic   [   0:0] snapshots$000$set_in_$040;
  logic   [   0:0] snapshots$000$set_in_$041;
  logic   [   0:0] snapshots$000$set_in_$042;
  logic   [   0:0] snapshots$000$set_in_$043;
  logic   [   0:0] snapshots$000$set_in_$044;
  logic   [   0:0] snapshots$000$set_in_$045;
  logic   [   0:0] snapshots$000$set_in_$046;
  logic   [   0:0] snapshots$000$set_in_$047;
  logic   [   0:0] snapshots$000$set_in_$048;
  logic   [   0:0] snapshots$000$set_in_$049;
  logic   [   0:0] snapshots$000$set_in_$050;
  logic   [   0:0] snapshots$000$set_in_$051;
  logic   [   0:0] snapshots$000$set_in_$052;
  logic   [   0:0] snapshots$000$set_in_$053;
  logic   [   0:0] snapshots$000$set_in_$054;
  logic   [   0:0] snapshots$000$set_in_$055;
  logic   [   0:0] snapshots$000$set_in_$056;
  logic   [   0:0] snapshots$000$set_in_$057;
  logic   [   0:0] snapshots$000$set_in_$058;
  logic   [   0:0] snapshots$000$set_in_$059;
  logic   [   0:0] snapshots$000$set_in_$060;
  logic   [   0:0] snapshots$000$set_in_$061;
  logic   [   0:0] snapshots$000$set_in_$062;
  logic   [   0:0] snapshots$000$set_call;
  logic   [   0:0] snapshots$000$clk;
  logic   [   5:0] snapshots$000$write_addr$000;
  logic   [   0:0] snapshots$000$write_call$000;
  logic   [   0:0] snapshots$000$write_data$000;
  logic   [   0:0] snapshots$000$reset;
  logic   [   0:0] snapshots$000$dump_out$000;
  logic   [   0:0] snapshots$000$dump_out$001;
  logic   [   0:0] snapshots$000$dump_out$002;
  logic   [   0:0] snapshots$000$dump_out$003;
  logic   [   0:0] snapshots$000$dump_out$004;
  logic   [   0:0] snapshots$000$dump_out$005;
  logic   [   0:0] snapshots$000$dump_out$006;
  logic   [   0:0] snapshots$000$dump_out$007;
  logic   [   0:0] snapshots$000$dump_out$008;
  logic   [   0:0] snapshots$000$dump_out$009;
  logic   [   0:0] snapshots$000$dump_out$010;
  logic   [   0:0] snapshots$000$dump_out$011;
  logic   [   0:0] snapshots$000$dump_out$012;
  logic   [   0:0] snapshots$000$dump_out$013;
  logic   [   0:0] snapshots$000$dump_out$014;
  logic   [   0:0] snapshots$000$dump_out$015;
  logic   [   0:0] snapshots$000$dump_out$016;
  logic   [   0:0] snapshots$000$dump_out$017;
  logic   [   0:0] snapshots$000$dump_out$018;
  logic   [   0:0] snapshots$000$dump_out$019;
  logic   [   0:0] snapshots$000$dump_out$020;
  logic   [   0:0] snapshots$000$dump_out$021;
  logic   [   0:0] snapshots$000$dump_out$022;
  logic   [   0:0] snapshots$000$dump_out$023;
  logic   [   0:0] snapshots$000$dump_out$024;
  logic   [   0:0] snapshots$000$dump_out$025;
  logic   [   0:0] snapshots$000$dump_out$026;
  logic   [   0:0] snapshots$000$dump_out$027;
  logic   [   0:0] snapshots$000$dump_out$028;
  logic   [   0:0] snapshots$000$dump_out$029;
  logic   [   0:0] snapshots$000$dump_out$030;
  logic   [   0:0] snapshots$000$dump_out$031;
  logic   [   0:0] snapshots$000$dump_out$032;
  logic   [   0:0] snapshots$000$dump_out$033;
  logic   [   0:0] snapshots$000$dump_out$034;
  logic   [   0:0] snapshots$000$dump_out$035;
  logic   [   0:0] snapshots$000$dump_out$036;
  logic   [   0:0] snapshots$000$dump_out$037;
  logic   [   0:0] snapshots$000$dump_out$038;
  logic   [   0:0] snapshots$000$dump_out$039;
  logic   [   0:0] snapshots$000$dump_out$040;
  logic   [   0:0] snapshots$000$dump_out$041;
  logic   [   0:0] snapshots$000$dump_out$042;
  logic   [   0:0] snapshots$000$dump_out$043;
  logic   [   0:0] snapshots$000$dump_out$044;
  logic   [   0:0] snapshots$000$dump_out$045;
  logic   [   0:0] snapshots$000$dump_out$046;
  logic   [   0:0] snapshots$000$dump_out$047;
  logic   [   0:0] snapshots$000$dump_out$048;
  logic   [   0:0] snapshots$000$dump_out$049;
  logic   [   0:0] snapshots$000$dump_out$050;
  logic   [   0:0] snapshots$000$dump_out$051;
  logic   [   0:0] snapshots$000$dump_out$052;
  logic   [   0:0] snapshots$000$dump_out$053;
  logic   [   0:0] snapshots$000$dump_out$054;
  logic   [   0:0] snapshots$000$dump_out$055;
  logic   [   0:0] snapshots$000$dump_out$056;
  logic   [   0:0] snapshots$000$dump_out$057;
  logic   [   0:0] snapshots$000$dump_out$058;
  logic   [   0:0] snapshots$000$dump_out$059;
  logic   [   0:0] snapshots$000$dump_out$060;
  logic   [   0:0] snapshots$000$dump_out$061;
  logic   [   0:0] snapshots$000$dump_out$062;

  RegisterFile_0x764ec1b6bf9dc34b snapshots$000
  (
    .set_in_$000    ( snapshots$000$set_in_$000 ),
    .set_in_$001    ( snapshots$000$set_in_$001 ),
    .set_in_$002    ( snapshots$000$set_in_$002 ),
    .set_in_$003    ( snapshots$000$set_in_$003 ),
    .set_in_$004    ( snapshots$000$set_in_$004 ),
    .set_in_$005    ( snapshots$000$set_in_$005 ),
    .set_in_$006    ( snapshots$000$set_in_$006 ),
    .set_in_$007    ( snapshots$000$set_in_$007 ),
    .set_in_$008    ( snapshots$000$set_in_$008 ),
    .set_in_$009    ( snapshots$000$set_in_$009 ),
    .set_in_$010    ( snapshots$000$set_in_$010 ),
    .set_in_$011    ( snapshots$000$set_in_$011 ),
    .set_in_$012    ( snapshots$000$set_in_$012 ),
    .set_in_$013    ( snapshots$000$set_in_$013 ),
    .set_in_$014    ( snapshots$000$set_in_$014 ),
    .set_in_$015    ( snapshots$000$set_in_$015 ),
    .set_in_$016    ( snapshots$000$set_in_$016 ),
    .set_in_$017    ( snapshots$000$set_in_$017 ),
    .set_in_$018    ( snapshots$000$set_in_$018 ),
    .set_in_$019    ( snapshots$000$set_in_$019 ),
    .set_in_$020    ( snapshots$000$set_in_$020 ),
    .set_in_$021    ( snapshots$000$set_in_$021 ),
    .set_in_$022    ( snapshots$000$set_in_$022 ),
    .set_in_$023    ( snapshots$000$set_in_$023 ),
    .set_in_$024    ( snapshots$000$set_in_$024 ),
    .set_in_$025    ( snapshots$000$set_in_$025 ),
    .set_in_$026    ( snapshots$000$set_in_$026 ),
    .set_in_$027    ( snapshots$000$set_in_$027 ),
    .set_in_$028    ( snapshots$000$set_in_$028 ),
    .set_in_$029    ( snapshots$000$set_in_$029 ),
    .set_in_$030    ( snapshots$000$set_in_$030 ),
    .set_in_$031    ( snapshots$000$set_in_$031 ),
    .set_in_$032    ( snapshots$000$set_in_$032 ),
    .set_in_$033    ( snapshots$000$set_in_$033 ),
    .set_in_$034    ( snapshots$000$set_in_$034 ),
    .set_in_$035    ( snapshots$000$set_in_$035 ),
    .set_in_$036    ( snapshots$000$set_in_$036 ),
    .set_in_$037    ( snapshots$000$set_in_$037 ),
    .set_in_$038    ( snapshots$000$set_in_$038 ),
    .set_in_$039    ( snapshots$000$set_in_$039 ),
    .set_in_$040    ( snapshots$000$set_in_$040 ),
    .set_in_$041    ( snapshots$000$set_in_$041 ),
    .set_in_$042    ( snapshots$000$set_in_$042 ),
    .set_in_$043    ( snapshots$000$set_in_$043 ),
    .set_in_$044    ( snapshots$000$set_in_$044 ),
    .set_in_$045    ( snapshots$000$set_in_$045 ),
    .set_in_$046    ( snapshots$000$set_in_$046 ),
    .set_in_$047    ( snapshots$000$set_in_$047 ),
    .set_in_$048    ( snapshots$000$set_in_$048 ),
    .set_in_$049    ( snapshots$000$set_in_$049 ),
    .set_in_$050    ( snapshots$000$set_in_$050 ),
    .set_in_$051    ( snapshots$000$set_in_$051 ),
    .set_in_$052    ( snapshots$000$set_in_$052 ),
    .set_in_$053    ( snapshots$000$set_in_$053 ),
    .set_in_$054    ( snapshots$000$set_in_$054 ),
    .set_in_$055    ( snapshots$000$set_in_$055 ),
    .set_in_$056    ( snapshots$000$set_in_$056 ),
    .set_in_$057    ( snapshots$000$set_in_$057 ),
    .set_in_$058    ( snapshots$000$set_in_$058 ),
    .set_in_$059    ( snapshots$000$set_in_$059 ),
    .set_in_$060    ( snapshots$000$set_in_$060 ),
    .set_in_$061    ( snapshots$000$set_in_$061 ),
    .set_in_$062    ( snapshots$000$set_in_$062 ),
    .set_call       ( snapshots$000$set_call ),
    .clk            ( snapshots$000$clk ),
    .write_addr$000 ( snapshots$000$write_addr$000 ),
    .write_call$000 ( snapshots$000$write_call$000 ),
    .write_data$000 ( snapshots$000$write_data$000 ),
    .reset          ( snapshots$000$reset ),
    .dump_out$000   ( snapshots$000$dump_out$000 ),
    .dump_out$001   ( snapshots$000$dump_out$001 ),
    .dump_out$002   ( snapshots$000$dump_out$002 ),
    .dump_out$003   ( snapshots$000$dump_out$003 ),
    .dump_out$004   ( snapshots$000$dump_out$004 ),
    .dump_out$005   ( snapshots$000$dump_out$005 ),
    .dump_out$006   ( snapshots$000$dump_out$006 ),
    .dump_out$007   ( snapshots$000$dump_out$007 ),
    .dump_out$008   ( snapshots$000$dump_out$008 ),
    .dump_out$009   ( snapshots$000$dump_out$009 ),
    .dump_out$010   ( snapshots$000$dump_out$010 ),
    .dump_out$011   ( snapshots$000$dump_out$011 ),
    .dump_out$012   ( snapshots$000$dump_out$012 ),
    .dump_out$013   ( snapshots$000$dump_out$013 ),
    .dump_out$014   ( snapshots$000$dump_out$014 ),
    .dump_out$015   ( snapshots$000$dump_out$015 ),
    .dump_out$016   ( snapshots$000$dump_out$016 ),
    .dump_out$017   ( snapshots$000$dump_out$017 ),
    .dump_out$018   ( snapshots$000$dump_out$018 ),
    .dump_out$019   ( snapshots$000$dump_out$019 ),
    .dump_out$020   ( snapshots$000$dump_out$020 ),
    .dump_out$021   ( snapshots$000$dump_out$021 ),
    .dump_out$022   ( snapshots$000$dump_out$022 ),
    .dump_out$023   ( snapshots$000$dump_out$023 ),
    .dump_out$024   ( snapshots$000$dump_out$024 ),
    .dump_out$025   ( snapshots$000$dump_out$025 ),
    .dump_out$026   ( snapshots$000$dump_out$026 ),
    .dump_out$027   ( snapshots$000$dump_out$027 ),
    .dump_out$028   ( snapshots$000$dump_out$028 ),
    .dump_out$029   ( snapshots$000$dump_out$029 ),
    .dump_out$030   ( snapshots$000$dump_out$030 ),
    .dump_out$031   ( snapshots$000$dump_out$031 ),
    .dump_out$032   ( snapshots$000$dump_out$032 ),
    .dump_out$033   ( snapshots$000$dump_out$033 ),
    .dump_out$034   ( snapshots$000$dump_out$034 ),
    .dump_out$035   ( snapshots$000$dump_out$035 ),
    .dump_out$036   ( snapshots$000$dump_out$036 ),
    .dump_out$037   ( snapshots$000$dump_out$037 ),
    .dump_out$038   ( snapshots$000$dump_out$038 ),
    .dump_out$039   ( snapshots$000$dump_out$039 ),
    .dump_out$040   ( snapshots$000$dump_out$040 ),
    .dump_out$041   ( snapshots$000$dump_out$041 ),
    .dump_out$042   ( snapshots$000$dump_out$042 ),
    .dump_out$043   ( snapshots$000$dump_out$043 ),
    .dump_out$044   ( snapshots$000$dump_out$044 ),
    .dump_out$045   ( snapshots$000$dump_out$045 ),
    .dump_out$046   ( snapshots$000$dump_out$046 ),
    .dump_out$047   ( snapshots$000$dump_out$047 ),
    .dump_out$048   ( snapshots$000$dump_out$048 ),
    .dump_out$049   ( snapshots$000$dump_out$049 ),
    .dump_out$050   ( snapshots$000$dump_out$050 ),
    .dump_out$051   ( snapshots$000$dump_out$051 ),
    .dump_out$052   ( snapshots$000$dump_out$052 ),
    .dump_out$053   ( snapshots$000$dump_out$053 ),
    .dump_out$054   ( snapshots$000$dump_out$054 ),
    .dump_out$055   ( snapshots$000$dump_out$055 ),
    .dump_out$056   ( snapshots$000$dump_out$056 ),
    .dump_out$057   ( snapshots$000$dump_out$057 ),
    .dump_out$058   ( snapshots$000$dump_out$058 ),
    .dump_out$059   ( snapshots$000$dump_out$059 ),
    .dump_out$060   ( snapshots$000$dump_out$060 ),
    .dump_out$061   ( snapshots$000$dump_out$061 ),
    .dump_out$062   ( snapshots$000$dump_out$062 )
  );

  // snapshots$001 temporaries
  logic   [   0:0] snapshots$001$set_in_$000;
  logic   [   0:0] snapshots$001$set_in_$001;
  logic   [   0:0] snapshots$001$set_in_$002;
  logic   [   0:0] snapshots$001$set_in_$003;
  logic   [   0:0] snapshots$001$set_in_$004;
  logic   [   0:0] snapshots$001$set_in_$005;
  logic   [   0:0] snapshots$001$set_in_$006;
  logic   [   0:0] snapshots$001$set_in_$007;
  logic   [   0:0] snapshots$001$set_in_$008;
  logic   [   0:0] snapshots$001$set_in_$009;
  logic   [   0:0] snapshots$001$set_in_$010;
  logic   [   0:0] snapshots$001$set_in_$011;
  logic   [   0:0] snapshots$001$set_in_$012;
  logic   [   0:0] snapshots$001$set_in_$013;
  logic   [   0:0] snapshots$001$set_in_$014;
  logic   [   0:0] snapshots$001$set_in_$015;
  logic   [   0:0] snapshots$001$set_in_$016;
  logic   [   0:0] snapshots$001$set_in_$017;
  logic   [   0:0] snapshots$001$set_in_$018;
  logic   [   0:0] snapshots$001$set_in_$019;
  logic   [   0:0] snapshots$001$set_in_$020;
  logic   [   0:0] snapshots$001$set_in_$021;
  logic   [   0:0] snapshots$001$set_in_$022;
  logic   [   0:0] snapshots$001$set_in_$023;
  logic   [   0:0] snapshots$001$set_in_$024;
  logic   [   0:0] snapshots$001$set_in_$025;
  logic   [   0:0] snapshots$001$set_in_$026;
  logic   [   0:0] snapshots$001$set_in_$027;
  logic   [   0:0] snapshots$001$set_in_$028;
  logic   [   0:0] snapshots$001$set_in_$029;
  logic   [   0:0] snapshots$001$set_in_$030;
  logic   [   0:0] snapshots$001$set_in_$031;
  logic   [   0:0] snapshots$001$set_in_$032;
  logic   [   0:0] snapshots$001$set_in_$033;
  logic   [   0:0] snapshots$001$set_in_$034;
  logic   [   0:0] snapshots$001$set_in_$035;
  logic   [   0:0] snapshots$001$set_in_$036;
  logic   [   0:0] snapshots$001$set_in_$037;
  logic   [   0:0] snapshots$001$set_in_$038;
  logic   [   0:0] snapshots$001$set_in_$039;
  logic   [   0:0] snapshots$001$set_in_$040;
  logic   [   0:0] snapshots$001$set_in_$041;
  logic   [   0:0] snapshots$001$set_in_$042;
  logic   [   0:0] snapshots$001$set_in_$043;
  logic   [   0:0] snapshots$001$set_in_$044;
  logic   [   0:0] snapshots$001$set_in_$045;
  logic   [   0:0] snapshots$001$set_in_$046;
  logic   [   0:0] snapshots$001$set_in_$047;
  logic   [   0:0] snapshots$001$set_in_$048;
  logic   [   0:0] snapshots$001$set_in_$049;
  logic   [   0:0] snapshots$001$set_in_$050;
  logic   [   0:0] snapshots$001$set_in_$051;
  logic   [   0:0] snapshots$001$set_in_$052;
  logic   [   0:0] snapshots$001$set_in_$053;
  logic   [   0:0] snapshots$001$set_in_$054;
  logic   [   0:0] snapshots$001$set_in_$055;
  logic   [   0:0] snapshots$001$set_in_$056;
  logic   [   0:0] snapshots$001$set_in_$057;
  logic   [   0:0] snapshots$001$set_in_$058;
  logic   [   0:0] snapshots$001$set_in_$059;
  logic   [   0:0] snapshots$001$set_in_$060;
  logic   [   0:0] snapshots$001$set_in_$061;
  logic   [   0:0] snapshots$001$set_in_$062;
  logic   [   0:0] snapshots$001$set_call;
  logic   [   0:0] snapshots$001$clk;
  logic   [   5:0] snapshots$001$write_addr$000;
  logic   [   0:0] snapshots$001$write_call$000;
  logic   [   0:0] snapshots$001$write_data$000;
  logic   [   0:0] snapshots$001$reset;
  logic   [   0:0] snapshots$001$dump_out$000;
  logic   [   0:0] snapshots$001$dump_out$001;
  logic   [   0:0] snapshots$001$dump_out$002;
  logic   [   0:0] snapshots$001$dump_out$003;
  logic   [   0:0] snapshots$001$dump_out$004;
  logic   [   0:0] snapshots$001$dump_out$005;
  logic   [   0:0] snapshots$001$dump_out$006;
  logic   [   0:0] snapshots$001$dump_out$007;
  logic   [   0:0] snapshots$001$dump_out$008;
  logic   [   0:0] snapshots$001$dump_out$009;
  logic   [   0:0] snapshots$001$dump_out$010;
  logic   [   0:0] snapshots$001$dump_out$011;
  logic   [   0:0] snapshots$001$dump_out$012;
  logic   [   0:0] snapshots$001$dump_out$013;
  logic   [   0:0] snapshots$001$dump_out$014;
  logic   [   0:0] snapshots$001$dump_out$015;
  logic   [   0:0] snapshots$001$dump_out$016;
  logic   [   0:0] snapshots$001$dump_out$017;
  logic   [   0:0] snapshots$001$dump_out$018;
  logic   [   0:0] snapshots$001$dump_out$019;
  logic   [   0:0] snapshots$001$dump_out$020;
  logic   [   0:0] snapshots$001$dump_out$021;
  logic   [   0:0] snapshots$001$dump_out$022;
  logic   [   0:0] snapshots$001$dump_out$023;
  logic   [   0:0] snapshots$001$dump_out$024;
  logic   [   0:0] snapshots$001$dump_out$025;
  logic   [   0:0] snapshots$001$dump_out$026;
  logic   [   0:0] snapshots$001$dump_out$027;
  logic   [   0:0] snapshots$001$dump_out$028;
  logic   [   0:0] snapshots$001$dump_out$029;
  logic   [   0:0] snapshots$001$dump_out$030;
  logic   [   0:0] snapshots$001$dump_out$031;
  logic   [   0:0] snapshots$001$dump_out$032;
  logic   [   0:0] snapshots$001$dump_out$033;
  logic   [   0:0] snapshots$001$dump_out$034;
  logic   [   0:0] snapshots$001$dump_out$035;
  logic   [   0:0] snapshots$001$dump_out$036;
  logic   [   0:0] snapshots$001$dump_out$037;
  logic   [   0:0] snapshots$001$dump_out$038;
  logic   [   0:0] snapshots$001$dump_out$039;
  logic   [   0:0] snapshots$001$dump_out$040;
  logic   [   0:0] snapshots$001$dump_out$041;
  logic   [   0:0] snapshots$001$dump_out$042;
  logic   [   0:0] snapshots$001$dump_out$043;
  logic   [   0:0] snapshots$001$dump_out$044;
  logic   [   0:0] snapshots$001$dump_out$045;
  logic   [   0:0] snapshots$001$dump_out$046;
  logic   [   0:0] snapshots$001$dump_out$047;
  logic   [   0:0] snapshots$001$dump_out$048;
  logic   [   0:0] snapshots$001$dump_out$049;
  logic   [   0:0] snapshots$001$dump_out$050;
  logic   [   0:0] snapshots$001$dump_out$051;
  logic   [   0:0] snapshots$001$dump_out$052;
  logic   [   0:0] snapshots$001$dump_out$053;
  logic   [   0:0] snapshots$001$dump_out$054;
  logic   [   0:0] snapshots$001$dump_out$055;
  logic   [   0:0] snapshots$001$dump_out$056;
  logic   [   0:0] snapshots$001$dump_out$057;
  logic   [   0:0] snapshots$001$dump_out$058;
  logic   [   0:0] snapshots$001$dump_out$059;
  logic   [   0:0] snapshots$001$dump_out$060;
  logic   [   0:0] snapshots$001$dump_out$061;
  logic   [   0:0] snapshots$001$dump_out$062;

  RegisterFile_0x764ec1b6bf9dc34b snapshots$001
  (
    .set_in_$000    ( snapshots$001$set_in_$000 ),
    .set_in_$001    ( snapshots$001$set_in_$001 ),
    .set_in_$002    ( snapshots$001$set_in_$002 ),
    .set_in_$003    ( snapshots$001$set_in_$003 ),
    .set_in_$004    ( snapshots$001$set_in_$004 ),
    .set_in_$005    ( snapshots$001$set_in_$005 ),
    .set_in_$006    ( snapshots$001$set_in_$006 ),
    .set_in_$007    ( snapshots$001$set_in_$007 ),
    .set_in_$008    ( snapshots$001$set_in_$008 ),
    .set_in_$009    ( snapshots$001$set_in_$009 ),
    .set_in_$010    ( snapshots$001$set_in_$010 ),
    .set_in_$011    ( snapshots$001$set_in_$011 ),
    .set_in_$012    ( snapshots$001$set_in_$012 ),
    .set_in_$013    ( snapshots$001$set_in_$013 ),
    .set_in_$014    ( snapshots$001$set_in_$014 ),
    .set_in_$015    ( snapshots$001$set_in_$015 ),
    .set_in_$016    ( snapshots$001$set_in_$016 ),
    .set_in_$017    ( snapshots$001$set_in_$017 ),
    .set_in_$018    ( snapshots$001$set_in_$018 ),
    .set_in_$019    ( snapshots$001$set_in_$019 ),
    .set_in_$020    ( snapshots$001$set_in_$020 ),
    .set_in_$021    ( snapshots$001$set_in_$021 ),
    .set_in_$022    ( snapshots$001$set_in_$022 ),
    .set_in_$023    ( snapshots$001$set_in_$023 ),
    .set_in_$024    ( snapshots$001$set_in_$024 ),
    .set_in_$025    ( snapshots$001$set_in_$025 ),
    .set_in_$026    ( snapshots$001$set_in_$026 ),
    .set_in_$027    ( snapshots$001$set_in_$027 ),
    .set_in_$028    ( snapshots$001$set_in_$028 ),
    .set_in_$029    ( snapshots$001$set_in_$029 ),
    .set_in_$030    ( snapshots$001$set_in_$030 ),
    .set_in_$031    ( snapshots$001$set_in_$031 ),
    .set_in_$032    ( snapshots$001$set_in_$032 ),
    .set_in_$033    ( snapshots$001$set_in_$033 ),
    .set_in_$034    ( snapshots$001$set_in_$034 ),
    .set_in_$035    ( snapshots$001$set_in_$035 ),
    .set_in_$036    ( snapshots$001$set_in_$036 ),
    .set_in_$037    ( snapshots$001$set_in_$037 ),
    .set_in_$038    ( snapshots$001$set_in_$038 ),
    .set_in_$039    ( snapshots$001$set_in_$039 ),
    .set_in_$040    ( snapshots$001$set_in_$040 ),
    .set_in_$041    ( snapshots$001$set_in_$041 ),
    .set_in_$042    ( snapshots$001$set_in_$042 ),
    .set_in_$043    ( snapshots$001$set_in_$043 ),
    .set_in_$044    ( snapshots$001$set_in_$044 ),
    .set_in_$045    ( snapshots$001$set_in_$045 ),
    .set_in_$046    ( snapshots$001$set_in_$046 ),
    .set_in_$047    ( snapshots$001$set_in_$047 ),
    .set_in_$048    ( snapshots$001$set_in_$048 ),
    .set_in_$049    ( snapshots$001$set_in_$049 ),
    .set_in_$050    ( snapshots$001$set_in_$050 ),
    .set_in_$051    ( snapshots$001$set_in_$051 ),
    .set_in_$052    ( snapshots$001$set_in_$052 ),
    .set_in_$053    ( snapshots$001$set_in_$053 ),
    .set_in_$054    ( snapshots$001$set_in_$054 ),
    .set_in_$055    ( snapshots$001$set_in_$055 ),
    .set_in_$056    ( snapshots$001$set_in_$056 ),
    .set_in_$057    ( snapshots$001$set_in_$057 ),
    .set_in_$058    ( snapshots$001$set_in_$058 ),
    .set_in_$059    ( snapshots$001$set_in_$059 ),
    .set_in_$060    ( snapshots$001$set_in_$060 ),
    .set_in_$061    ( snapshots$001$set_in_$061 ),
    .set_in_$062    ( snapshots$001$set_in_$062 ),
    .set_call       ( snapshots$001$set_call ),
    .clk            ( snapshots$001$clk ),
    .write_addr$000 ( snapshots$001$write_addr$000 ),
    .write_call$000 ( snapshots$001$write_call$000 ),
    .write_data$000 ( snapshots$001$write_data$000 ),
    .reset          ( snapshots$001$reset ),
    .dump_out$000   ( snapshots$001$dump_out$000 ),
    .dump_out$001   ( snapshots$001$dump_out$001 ),
    .dump_out$002   ( snapshots$001$dump_out$002 ),
    .dump_out$003   ( snapshots$001$dump_out$003 ),
    .dump_out$004   ( snapshots$001$dump_out$004 ),
    .dump_out$005   ( snapshots$001$dump_out$005 ),
    .dump_out$006   ( snapshots$001$dump_out$006 ),
    .dump_out$007   ( snapshots$001$dump_out$007 ),
    .dump_out$008   ( snapshots$001$dump_out$008 ),
    .dump_out$009   ( snapshots$001$dump_out$009 ),
    .dump_out$010   ( snapshots$001$dump_out$010 ),
    .dump_out$011   ( snapshots$001$dump_out$011 ),
    .dump_out$012   ( snapshots$001$dump_out$012 ),
    .dump_out$013   ( snapshots$001$dump_out$013 ),
    .dump_out$014   ( snapshots$001$dump_out$014 ),
    .dump_out$015   ( snapshots$001$dump_out$015 ),
    .dump_out$016   ( snapshots$001$dump_out$016 ),
    .dump_out$017   ( snapshots$001$dump_out$017 ),
    .dump_out$018   ( snapshots$001$dump_out$018 ),
    .dump_out$019   ( snapshots$001$dump_out$019 ),
    .dump_out$020   ( snapshots$001$dump_out$020 ),
    .dump_out$021   ( snapshots$001$dump_out$021 ),
    .dump_out$022   ( snapshots$001$dump_out$022 ),
    .dump_out$023   ( snapshots$001$dump_out$023 ),
    .dump_out$024   ( snapshots$001$dump_out$024 ),
    .dump_out$025   ( snapshots$001$dump_out$025 ),
    .dump_out$026   ( snapshots$001$dump_out$026 ),
    .dump_out$027   ( snapshots$001$dump_out$027 ),
    .dump_out$028   ( snapshots$001$dump_out$028 ),
    .dump_out$029   ( snapshots$001$dump_out$029 ),
    .dump_out$030   ( snapshots$001$dump_out$030 ),
    .dump_out$031   ( snapshots$001$dump_out$031 ),
    .dump_out$032   ( snapshots$001$dump_out$032 ),
    .dump_out$033   ( snapshots$001$dump_out$033 ),
    .dump_out$034   ( snapshots$001$dump_out$034 ),
    .dump_out$035   ( snapshots$001$dump_out$035 ),
    .dump_out$036   ( snapshots$001$dump_out$036 ),
    .dump_out$037   ( snapshots$001$dump_out$037 ),
    .dump_out$038   ( snapshots$001$dump_out$038 ),
    .dump_out$039   ( snapshots$001$dump_out$039 ),
    .dump_out$040   ( snapshots$001$dump_out$040 ),
    .dump_out$041   ( snapshots$001$dump_out$041 ),
    .dump_out$042   ( snapshots$001$dump_out$042 ),
    .dump_out$043   ( snapshots$001$dump_out$043 ),
    .dump_out$044   ( snapshots$001$dump_out$044 ),
    .dump_out$045   ( snapshots$001$dump_out$045 ),
    .dump_out$046   ( snapshots$001$dump_out$046 ),
    .dump_out$047   ( snapshots$001$dump_out$047 ),
    .dump_out$048   ( snapshots$001$dump_out$048 ),
    .dump_out$049   ( snapshots$001$dump_out$049 ),
    .dump_out$050   ( snapshots$001$dump_out$050 ),
    .dump_out$051   ( snapshots$001$dump_out$051 ),
    .dump_out$052   ( snapshots$001$dump_out$052 ),
    .dump_out$053   ( snapshots$001$dump_out$053 ),
    .dump_out$054   ( snapshots$001$dump_out$054 ),
    .dump_out$055   ( snapshots$001$dump_out$055 ),
    .dump_out$056   ( snapshots$001$dump_out$056 ),
    .dump_out$057   ( snapshots$001$dump_out$057 ),
    .dump_out$058   ( snapshots$001$dump_out$058 ),
    .dump_out$059   ( snapshots$001$dump_out$059 ),
    .dump_out$060   ( snapshots$001$dump_out$060 ),
    .dump_out$061   ( snapshots$001$dump_out$061 ),
    .dump_out$062   ( snapshots$001$dump_out$062 )
  );

  // dump_mux temporaries
  logic   [  62:0] dump_mux$mux_in_$000;
  logic   [  62:0] dump_mux$mux_in_$001;
  logic   [   0:0] dump_mux$clk;
  logic   [   0:0] dump_mux$reset;
  logic   [   0:0] dump_mux$mux_select;
  logic   [  62:0] dump_mux$mux_out;

  Mux_0x7af68b5383bacfb2 dump_mux
  (
    .mux_in_$000 ( dump_mux$mux_in_$000 ),
    .mux_in_$001 ( dump_mux$mux_in_$001 ),
    .clk         ( dump_mux$clk ),
    .reset       ( dump_mux$reset ),
    .mux_select  ( dump_mux$mux_select ),
    .mux_out     ( dump_mux$mux_out )
  );

  // free_list temporaries
  logic   [  62:0] free_list$set_state;
  logic   [   0:0] free_list$clk;
  logic   [   0:0] free_list$free_call$000;
  logic   [   0:0] free_list$free_call$001;
  logic   [  62:0] free_list$release_mask;
  logic   [   0:0] free_list$alloc_call$000;
  logic   [   0:0] free_list$reset;
  logic   [   0:0] free_list$set_call;
  logic   [   5:0] free_list$free_index$000;
  logic   [   5:0] free_list$free_index$001;
  logic   [  62:0] free_list$alloc_mask$000;
  logic   [   0:0] free_list$alloc_rdy$000;
  logic   [   5:0] free_list$alloc_index$000;

  FreeList_0x2dd76b08b1ccb6ed free_list
  (
    .set_state       ( free_list$set_state ),
    .release_call    ( free_list$release_call ),
    .clk             ( free_list$clk ),
    .free_call$000   ( free_list$free_call$000 ),
    .free_call$001   ( free_list$free_call$001 ),
    .release_mask    ( free_list$release_mask ),
    .alloc_call$000  ( free_list$alloc_call$000 ),
    .reset           ( free_list$reset ),
    .set_call        ( free_list$set_call ),
    .free_index$000  ( free_list$free_index$000 ),
    .free_index$001  ( free_list$free_index$001 ),
    .alloc_mask$000  ( free_list$alloc_mask$000 ),
    .alloc_rdy$000   ( free_list$alloc_rdy$000 ),
    .alloc_index$000 ( free_list$alloc_index$000 )
  );

  // snapshot_packers$000 temporaries
  logic   [   0:0] snapshot_packers$000$clk;
  logic   [   0:0] snapshot_packers$000$pack_in_$000;
  logic   [   0:0] snapshot_packers$000$pack_in_$001;
  logic   [   0:0] snapshot_packers$000$pack_in_$002;
  logic   [   0:0] snapshot_packers$000$pack_in_$003;
  logic   [   0:0] snapshot_packers$000$pack_in_$004;
  logic   [   0:0] snapshot_packers$000$pack_in_$005;
  logic   [   0:0] snapshot_packers$000$pack_in_$006;
  logic   [   0:0] snapshot_packers$000$pack_in_$007;
  logic   [   0:0] snapshot_packers$000$pack_in_$008;
  logic   [   0:0] snapshot_packers$000$pack_in_$009;
  logic   [   0:0] snapshot_packers$000$pack_in_$010;
  logic   [   0:0] snapshot_packers$000$pack_in_$011;
  logic   [   0:0] snapshot_packers$000$pack_in_$012;
  logic   [   0:0] snapshot_packers$000$pack_in_$013;
  logic   [   0:0] snapshot_packers$000$pack_in_$014;
  logic   [   0:0] snapshot_packers$000$pack_in_$015;
  logic   [   0:0] snapshot_packers$000$pack_in_$016;
  logic   [   0:0] snapshot_packers$000$pack_in_$017;
  logic   [   0:0] snapshot_packers$000$pack_in_$018;
  logic   [   0:0] snapshot_packers$000$pack_in_$019;
  logic   [   0:0] snapshot_packers$000$pack_in_$020;
  logic   [   0:0] snapshot_packers$000$pack_in_$021;
  logic   [   0:0] snapshot_packers$000$pack_in_$022;
  logic   [   0:0] snapshot_packers$000$pack_in_$023;
  logic   [   0:0] snapshot_packers$000$pack_in_$024;
  logic   [   0:0] snapshot_packers$000$pack_in_$025;
  logic   [   0:0] snapshot_packers$000$pack_in_$026;
  logic   [   0:0] snapshot_packers$000$pack_in_$027;
  logic   [   0:0] snapshot_packers$000$pack_in_$028;
  logic   [   0:0] snapshot_packers$000$pack_in_$029;
  logic   [   0:0] snapshot_packers$000$pack_in_$030;
  logic   [   0:0] snapshot_packers$000$pack_in_$031;
  logic   [   0:0] snapshot_packers$000$pack_in_$032;
  logic   [   0:0] snapshot_packers$000$pack_in_$033;
  logic   [   0:0] snapshot_packers$000$pack_in_$034;
  logic   [   0:0] snapshot_packers$000$pack_in_$035;
  logic   [   0:0] snapshot_packers$000$pack_in_$036;
  logic   [   0:0] snapshot_packers$000$pack_in_$037;
  logic   [   0:0] snapshot_packers$000$pack_in_$038;
  logic   [   0:0] snapshot_packers$000$pack_in_$039;
  logic   [   0:0] snapshot_packers$000$pack_in_$040;
  logic   [   0:0] snapshot_packers$000$pack_in_$041;
  logic   [   0:0] snapshot_packers$000$pack_in_$042;
  logic   [   0:0] snapshot_packers$000$pack_in_$043;
  logic   [   0:0] snapshot_packers$000$pack_in_$044;
  logic   [   0:0] snapshot_packers$000$pack_in_$045;
  logic   [   0:0] snapshot_packers$000$pack_in_$046;
  logic   [   0:0] snapshot_packers$000$pack_in_$047;
  logic   [   0:0] snapshot_packers$000$pack_in_$048;
  logic   [   0:0] snapshot_packers$000$pack_in_$049;
  logic   [   0:0] snapshot_packers$000$pack_in_$050;
  logic   [   0:0] snapshot_packers$000$pack_in_$051;
  logic   [   0:0] snapshot_packers$000$pack_in_$052;
  logic   [   0:0] snapshot_packers$000$pack_in_$053;
  logic   [   0:0] snapshot_packers$000$pack_in_$054;
  logic   [   0:0] snapshot_packers$000$pack_in_$055;
  logic   [   0:0] snapshot_packers$000$pack_in_$056;
  logic   [   0:0] snapshot_packers$000$pack_in_$057;
  logic   [   0:0] snapshot_packers$000$pack_in_$058;
  logic   [   0:0] snapshot_packers$000$pack_in_$059;
  logic   [   0:0] snapshot_packers$000$pack_in_$060;
  logic   [   0:0] snapshot_packers$000$pack_in_$061;
  logic   [   0:0] snapshot_packers$000$pack_in_$062;
  logic   [   0:0] snapshot_packers$000$reset;
  logic   [  62:0] snapshot_packers$000$pack_packed;

  Packer_0x5417ceb8bd59f204 snapshot_packers$000
  (
    .clk          ( snapshot_packers$000$clk ),
    .pack_in_$000 ( snapshot_packers$000$pack_in_$000 ),
    .pack_in_$001 ( snapshot_packers$000$pack_in_$001 ),
    .pack_in_$002 ( snapshot_packers$000$pack_in_$002 ),
    .pack_in_$003 ( snapshot_packers$000$pack_in_$003 ),
    .pack_in_$004 ( snapshot_packers$000$pack_in_$004 ),
    .pack_in_$005 ( snapshot_packers$000$pack_in_$005 ),
    .pack_in_$006 ( snapshot_packers$000$pack_in_$006 ),
    .pack_in_$007 ( snapshot_packers$000$pack_in_$007 ),
    .pack_in_$008 ( snapshot_packers$000$pack_in_$008 ),
    .pack_in_$009 ( snapshot_packers$000$pack_in_$009 ),
    .pack_in_$010 ( snapshot_packers$000$pack_in_$010 ),
    .pack_in_$011 ( snapshot_packers$000$pack_in_$011 ),
    .pack_in_$012 ( snapshot_packers$000$pack_in_$012 ),
    .pack_in_$013 ( snapshot_packers$000$pack_in_$013 ),
    .pack_in_$014 ( snapshot_packers$000$pack_in_$014 ),
    .pack_in_$015 ( snapshot_packers$000$pack_in_$015 ),
    .pack_in_$016 ( snapshot_packers$000$pack_in_$016 ),
    .pack_in_$017 ( snapshot_packers$000$pack_in_$017 ),
    .pack_in_$018 ( snapshot_packers$000$pack_in_$018 ),
    .pack_in_$019 ( snapshot_packers$000$pack_in_$019 ),
    .pack_in_$020 ( snapshot_packers$000$pack_in_$020 ),
    .pack_in_$021 ( snapshot_packers$000$pack_in_$021 ),
    .pack_in_$022 ( snapshot_packers$000$pack_in_$022 ),
    .pack_in_$023 ( snapshot_packers$000$pack_in_$023 ),
    .pack_in_$024 ( snapshot_packers$000$pack_in_$024 ),
    .pack_in_$025 ( snapshot_packers$000$pack_in_$025 ),
    .pack_in_$026 ( snapshot_packers$000$pack_in_$026 ),
    .pack_in_$027 ( snapshot_packers$000$pack_in_$027 ),
    .pack_in_$028 ( snapshot_packers$000$pack_in_$028 ),
    .pack_in_$029 ( snapshot_packers$000$pack_in_$029 ),
    .pack_in_$030 ( snapshot_packers$000$pack_in_$030 ),
    .pack_in_$031 ( snapshot_packers$000$pack_in_$031 ),
    .pack_in_$032 ( snapshot_packers$000$pack_in_$032 ),
    .pack_in_$033 ( snapshot_packers$000$pack_in_$033 ),
    .pack_in_$034 ( snapshot_packers$000$pack_in_$034 ),
    .pack_in_$035 ( snapshot_packers$000$pack_in_$035 ),
    .pack_in_$036 ( snapshot_packers$000$pack_in_$036 ),
    .pack_in_$037 ( snapshot_packers$000$pack_in_$037 ),
    .pack_in_$038 ( snapshot_packers$000$pack_in_$038 ),
    .pack_in_$039 ( snapshot_packers$000$pack_in_$039 ),
    .pack_in_$040 ( snapshot_packers$000$pack_in_$040 ),
    .pack_in_$041 ( snapshot_packers$000$pack_in_$041 ),
    .pack_in_$042 ( snapshot_packers$000$pack_in_$042 ),
    .pack_in_$043 ( snapshot_packers$000$pack_in_$043 ),
    .pack_in_$044 ( snapshot_packers$000$pack_in_$044 ),
    .pack_in_$045 ( snapshot_packers$000$pack_in_$045 ),
    .pack_in_$046 ( snapshot_packers$000$pack_in_$046 ),
    .pack_in_$047 ( snapshot_packers$000$pack_in_$047 ),
    .pack_in_$048 ( snapshot_packers$000$pack_in_$048 ),
    .pack_in_$049 ( snapshot_packers$000$pack_in_$049 ),
    .pack_in_$050 ( snapshot_packers$000$pack_in_$050 ),
    .pack_in_$051 ( snapshot_packers$000$pack_in_$051 ),
    .pack_in_$052 ( snapshot_packers$000$pack_in_$052 ),
    .pack_in_$053 ( snapshot_packers$000$pack_in_$053 ),
    .pack_in_$054 ( snapshot_packers$000$pack_in_$054 ),
    .pack_in_$055 ( snapshot_packers$000$pack_in_$055 ),
    .pack_in_$056 ( snapshot_packers$000$pack_in_$056 ),
    .pack_in_$057 ( snapshot_packers$000$pack_in_$057 ),
    .pack_in_$058 ( snapshot_packers$000$pack_in_$058 ),
    .pack_in_$059 ( snapshot_packers$000$pack_in_$059 ),
    .pack_in_$060 ( snapshot_packers$000$pack_in_$060 ),
    .pack_in_$061 ( snapshot_packers$000$pack_in_$061 ),
    .pack_in_$062 ( snapshot_packers$000$pack_in_$062 ),
    .reset        ( snapshot_packers$000$reset ),
    .pack_packed  ( snapshot_packers$000$pack_packed )
  );

  // snapshot_packers$001 temporaries
  logic   [   0:0] snapshot_packers$001$clk;
  logic   [   0:0] snapshot_packers$001$pack_in_$000;
  logic   [   0:0] snapshot_packers$001$pack_in_$001;
  logic   [   0:0] snapshot_packers$001$pack_in_$002;
  logic   [   0:0] snapshot_packers$001$pack_in_$003;
  logic   [   0:0] snapshot_packers$001$pack_in_$004;
  logic   [   0:0] snapshot_packers$001$pack_in_$005;
  logic   [   0:0] snapshot_packers$001$pack_in_$006;
  logic   [   0:0] snapshot_packers$001$pack_in_$007;
  logic   [   0:0] snapshot_packers$001$pack_in_$008;
  logic   [   0:0] snapshot_packers$001$pack_in_$009;
  logic   [   0:0] snapshot_packers$001$pack_in_$010;
  logic   [   0:0] snapshot_packers$001$pack_in_$011;
  logic   [   0:0] snapshot_packers$001$pack_in_$012;
  logic   [   0:0] snapshot_packers$001$pack_in_$013;
  logic   [   0:0] snapshot_packers$001$pack_in_$014;
  logic   [   0:0] snapshot_packers$001$pack_in_$015;
  logic   [   0:0] snapshot_packers$001$pack_in_$016;
  logic   [   0:0] snapshot_packers$001$pack_in_$017;
  logic   [   0:0] snapshot_packers$001$pack_in_$018;
  logic   [   0:0] snapshot_packers$001$pack_in_$019;
  logic   [   0:0] snapshot_packers$001$pack_in_$020;
  logic   [   0:0] snapshot_packers$001$pack_in_$021;
  logic   [   0:0] snapshot_packers$001$pack_in_$022;
  logic   [   0:0] snapshot_packers$001$pack_in_$023;
  logic   [   0:0] snapshot_packers$001$pack_in_$024;
  logic   [   0:0] snapshot_packers$001$pack_in_$025;
  logic   [   0:0] snapshot_packers$001$pack_in_$026;
  logic   [   0:0] snapshot_packers$001$pack_in_$027;
  logic   [   0:0] snapshot_packers$001$pack_in_$028;
  logic   [   0:0] snapshot_packers$001$pack_in_$029;
  logic   [   0:0] snapshot_packers$001$pack_in_$030;
  logic   [   0:0] snapshot_packers$001$pack_in_$031;
  logic   [   0:0] snapshot_packers$001$pack_in_$032;
  logic   [   0:0] snapshot_packers$001$pack_in_$033;
  logic   [   0:0] snapshot_packers$001$pack_in_$034;
  logic   [   0:0] snapshot_packers$001$pack_in_$035;
  logic   [   0:0] snapshot_packers$001$pack_in_$036;
  logic   [   0:0] snapshot_packers$001$pack_in_$037;
  logic   [   0:0] snapshot_packers$001$pack_in_$038;
  logic   [   0:0] snapshot_packers$001$pack_in_$039;
  logic   [   0:0] snapshot_packers$001$pack_in_$040;
  logic   [   0:0] snapshot_packers$001$pack_in_$041;
  logic   [   0:0] snapshot_packers$001$pack_in_$042;
  logic   [   0:0] snapshot_packers$001$pack_in_$043;
  logic   [   0:0] snapshot_packers$001$pack_in_$044;
  logic   [   0:0] snapshot_packers$001$pack_in_$045;
  logic   [   0:0] snapshot_packers$001$pack_in_$046;
  logic   [   0:0] snapshot_packers$001$pack_in_$047;
  logic   [   0:0] snapshot_packers$001$pack_in_$048;
  logic   [   0:0] snapshot_packers$001$pack_in_$049;
  logic   [   0:0] snapshot_packers$001$pack_in_$050;
  logic   [   0:0] snapshot_packers$001$pack_in_$051;
  logic   [   0:0] snapshot_packers$001$pack_in_$052;
  logic   [   0:0] snapshot_packers$001$pack_in_$053;
  logic   [   0:0] snapshot_packers$001$pack_in_$054;
  logic   [   0:0] snapshot_packers$001$pack_in_$055;
  logic   [   0:0] snapshot_packers$001$pack_in_$056;
  logic   [   0:0] snapshot_packers$001$pack_in_$057;
  logic   [   0:0] snapshot_packers$001$pack_in_$058;
  logic   [   0:0] snapshot_packers$001$pack_in_$059;
  logic   [   0:0] snapshot_packers$001$pack_in_$060;
  logic   [   0:0] snapshot_packers$001$pack_in_$061;
  logic   [   0:0] snapshot_packers$001$pack_in_$062;
  logic   [   0:0] snapshot_packers$001$reset;
  logic   [  62:0] snapshot_packers$001$pack_packed;

  Packer_0x5417ceb8bd59f204 snapshot_packers$001
  (
    .clk          ( snapshot_packers$001$clk ),
    .pack_in_$000 ( snapshot_packers$001$pack_in_$000 ),
    .pack_in_$001 ( snapshot_packers$001$pack_in_$001 ),
    .pack_in_$002 ( snapshot_packers$001$pack_in_$002 ),
    .pack_in_$003 ( snapshot_packers$001$pack_in_$003 ),
    .pack_in_$004 ( snapshot_packers$001$pack_in_$004 ),
    .pack_in_$005 ( snapshot_packers$001$pack_in_$005 ),
    .pack_in_$006 ( snapshot_packers$001$pack_in_$006 ),
    .pack_in_$007 ( snapshot_packers$001$pack_in_$007 ),
    .pack_in_$008 ( snapshot_packers$001$pack_in_$008 ),
    .pack_in_$009 ( snapshot_packers$001$pack_in_$009 ),
    .pack_in_$010 ( snapshot_packers$001$pack_in_$010 ),
    .pack_in_$011 ( snapshot_packers$001$pack_in_$011 ),
    .pack_in_$012 ( snapshot_packers$001$pack_in_$012 ),
    .pack_in_$013 ( snapshot_packers$001$pack_in_$013 ),
    .pack_in_$014 ( snapshot_packers$001$pack_in_$014 ),
    .pack_in_$015 ( snapshot_packers$001$pack_in_$015 ),
    .pack_in_$016 ( snapshot_packers$001$pack_in_$016 ),
    .pack_in_$017 ( snapshot_packers$001$pack_in_$017 ),
    .pack_in_$018 ( snapshot_packers$001$pack_in_$018 ),
    .pack_in_$019 ( snapshot_packers$001$pack_in_$019 ),
    .pack_in_$020 ( snapshot_packers$001$pack_in_$020 ),
    .pack_in_$021 ( snapshot_packers$001$pack_in_$021 ),
    .pack_in_$022 ( snapshot_packers$001$pack_in_$022 ),
    .pack_in_$023 ( snapshot_packers$001$pack_in_$023 ),
    .pack_in_$024 ( snapshot_packers$001$pack_in_$024 ),
    .pack_in_$025 ( snapshot_packers$001$pack_in_$025 ),
    .pack_in_$026 ( snapshot_packers$001$pack_in_$026 ),
    .pack_in_$027 ( snapshot_packers$001$pack_in_$027 ),
    .pack_in_$028 ( snapshot_packers$001$pack_in_$028 ),
    .pack_in_$029 ( snapshot_packers$001$pack_in_$029 ),
    .pack_in_$030 ( snapshot_packers$001$pack_in_$030 ),
    .pack_in_$031 ( snapshot_packers$001$pack_in_$031 ),
    .pack_in_$032 ( snapshot_packers$001$pack_in_$032 ),
    .pack_in_$033 ( snapshot_packers$001$pack_in_$033 ),
    .pack_in_$034 ( snapshot_packers$001$pack_in_$034 ),
    .pack_in_$035 ( snapshot_packers$001$pack_in_$035 ),
    .pack_in_$036 ( snapshot_packers$001$pack_in_$036 ),
    .pack_in_$037 ( snapshot_packers$001$pack_in_$037 ),
    .pack_in_$038 ( snapshot_packers$001$pack_in_$038 ),
    .pack_in_$039 ( snapshot_packers$001$pack_in_$039 ),
    .pack_in_$040 ( snapshot_packers$001$pack_in_$040 ),
    .pack_in_$041 ( snapshot_packers$001$pack_in_$041 ),
    .pack_in_$042 ( snapshot_packers$001$pack_in_$042 ),
    .pack_in_$043 ( snapshot_packers$001$pack_in_$043 ),
    .pack_in_$044 ( snapshot_packers$001$pack_in_$044 ),
    .pack_in_$045 ( snapshot_packers$001$pack_in_$045 ),
    .pack_in_$046 ( snapshot_packers$001$pack_in_$046 ),
    .pack_in_$047 ( snapshot_packers$001$pack_in_$047 ),
    .pack_in_$048 ( snapshot_packers$001$pack_in_$048 ),
    .pack_in_$049 ( snapshot_packers$001$pack_in_$049 ),
    .pack_in_$050 ( snapshot_packers$001$pack_in_$050 ),
    .pack_in_$051 ( snapshot_packers$001$pack_in_$051 ),
    .pack_in_$052 ( snapshot_packers$001$pack_in_$052 ),
    .pack_in_$053 ( snapshot_packers$001$pack_in_$053 ),
    .pack_in_$054 ( snapshot_packers$001$pack_in_$054 ),
    .pack_in_$055 ( snapshot_packers$001$pack_in_$055 ),
    .pack_in_$056 ( snapshot_packers$001$pack_in_$056 ),
    .pack_in_$057 ( snapshot_packers$001$pack_in_$057 ),
    .pack_in_$058 ( snapshot_packers$001$pack_in_$058 ),
    .pack_in_$059 ( snapshot_packers$001$pack_in_$059 ),
    .pack_in_$060 ( snapshot_packers$001$pack_in_$060 ),
    .pack_in_$061 ( snapshot_packers$001$pack_in_$061 ),
    .pack_in_$062 ( snapshot_packers$001$pack_in_$062 ),
    .reset        ( snapshot_packers$001$reset ),
    .pack_packed  ( snapshot_packers$001$pack_packed )
  );

  // clean_mux temporaries
  logic   [  62:0] clean_mux$mux_in_$000;
  logic   [  62:0] clean_mux$mux_in_$001;
  logic   [   0:0] clean_mux$clk;
  logic   [   0:0] clean_mux$reset;
  logic   [   0:0] clean_mux$mux_select;
  logic   [  62:0] clean_mux$mux_out;

  Mux_0x7af68b5383bacfb2 clean_mux
  (
    .mux_in_$000 ( clean_mux$mux_in_$000 ),
    .mux_in_$001 ( clean_mux$mux_in_$001 ),
    .clk         ( clean_mux$clk ),
    .reset       ( clean_mux$reset ),
    .mux_select  ( clean_mux$mux_select ),
    .mux_out     ( clean_mux$mux_out )
  );

  // signal connections
  assign alloc_index$000                   = free_list$alloc_index$000;
  assign alloc_mask$000                    = free_list$alloc_mask$000;
  assign alloc_rdy$000                     = free_list$alloc_rdy$000;
  assign clean_mux$clk                     = clk;
  assign clean_mux$reset                   = reset;
  assign dump_mux$clk                      = clk;
  assign dump_mux$mux_in_$000              = snapshot_packers$000$pack_packed;
  assign dump_mux$mux_in_$001              = snapshot_packers$001$pack_packed;
  assign dump_mux$mux_select               = revert_allocs_source_id;
  assign dump_mux$reset                    = reset;
  assign free_list$alloc_call$000          = alloc_call$000;
  assign free_list$clk                     = clk;
  assign free_list$free_call$000           = free_call$000;
  assign free_list$free_call$001           = free_call$001;
  assign free_list$free_index$000          = free_index$000;
  assign free_list$free_index$001          = free_index$001;
  assign free_list$release_mask            = dump_mux$mux_out;
  assign free_list$reset                   = reset;
  assign free_list$set_call                = set_call;
  assign free_list$set_state               = set_state;
  assign snapshot_packers$000$clk          = clk;
  assign snapshot_packers$000$pack_in_$000 = snapshots$000$dump_out$000;
  assign snapshot_packers$000$pack_in_$001 = snapshots$000$dump_out$001;
  assign snapshot_packers$000$pack_in_$002 = snapshots$000$dump_out$002;
  assign snapshot_packers$000$pack_in_$003 = snapshots$000$dump_out$003;
  assign snapshot_packers$000$pack_in_$004 = snapshots$000$dump_out$004;
  assign snapshot_packers$000$pack_in_$005 = snapshots$000$dump_out$005;
  assign snapshot_packers$000$pack_in_$006 = snapshots$000$dump_out$006;
  assign snapshot_packers$000$pack_in_$007 = snapshots$000$dump_out$007;
  assign snapshot_packers$000$pack_in_$008 = snapshots$000$dump_out$008;
  assign snapshot_packers$000$pack_in_$009 = snapshots$000$dump_out$009;
  assign snapshot_packers$000$pack_in_$010 = snapshots$000$dump_out$010;
  assign snapshot_packers$000$pack_in_$011 = snapshots$000$dump_out$011;
  assign snapshot_packers$000$pack_in_$012 = snapshots$000$dump_out$012;
  assign snapshot_packers$000$pack_in_$013 = snapshots$000$dump_out$013;
  assign snapshot_packers$000$pack_in_$014 = snapshots$000$dump_out$014;
  assign snapshot_packers$000$pack_in_$015 = snapshots$000$dump_out$015;
  assign snapshot_packers$000$pack_in_$016 = snapshots$000$dump_out$016;
  assign snapshot_packers$000$pack_in_$017 = snapshots$000$dump_out$017;
  assign snapshot_packers$000$pack_in_$018 = snapshots$000$dump_out$018;
  assign snapshot_packers$000$pack_in_$019 = snapshots$000$dump_out$019;
  assign snapshot_packers$000$pack_in_$020 = snapshots$000$dump_out$020;
  assign snapshot_packers$000$pack_in_$021 = snapshots$000$dump_out$021;
  assign snapshot_packers$000$pack_in_$022 = snapshots$000$dump_out$022;
  assign snapshot_packers$000$pack_in_$023 = snapshots$000$dump_out$023;
  assign snapshot_packers$000$pack_in_$024 = snapshots$000$dump_out$024;
  assign snapshot_packers$000$pack_in_$025 = snapshots$000$dump_out$025;
  assign snapshot_packers$000$pack_in_$026 = snapshots$000$dump_out$026;
  assign snapshot_packers$000$pack_in_$027 = snapshots$000$dump_out$027;
  assign snapshot_packers$000$pack_in_$028 = snapshots$000$dump_out$028;
  assign snapshot_packers$000$pack_in_$029 = snapshots$000$dump_out$029;
  assign snapshot_packers$000$pack_in_$030 = snapshots$000$dump_out$030;
  assign snapshot_packers$000$pack_in_$031 = snapshots$000$dump_out$031;
  assign snapshot_packers$000$pack_in_$032 = snapshots$000$dump_out$032;
  assign snapshot_packers$000$pack_in_$033 = snapshots$000$dump_out$033;
  assign snapshot_packers$000$pack_in_$034 = snapshots$000$dump_out$034;
  assign snapshot_packers$000$pack_in_$035 = snapshots$000$dump_out$035;
  assign snapshot_packers$000$pack_in_$036 = snapshots$000$dump_out$036;
  assign snapshot_packers$000$pack_in_$037 = snapshots$000$dump_out$037;
  assign snapshot_packers$000$pack_in_$038 = snapshots$000$dump_out$038;
  assign snapshot_packers$000$pack_in_$039 = snapshots$000$dump_out$039;
  assign snapshot_packers$000$pack_in_$040 = snapshots$000$dump_out$040;
  assign snapshot_packers$000$pack_in_$041 = snapshots$000$dump_out$041;
  assign snapshot_packers$000$pack_in_$042 = snapshots$000$dump_out$042;
  assign snapshot_packers$000$pack_in_$043 = snapshots$000$dump_out$043;
  assign snapshot_packers$000$pack_in_$044 = snapshots$000$dump_out$044;
  assign snapshot_packers$000$pack_in_$045 = snapshots$000$dump_out$045;
  assign snapshot_packers$000$pack_in_$046 = snapshots$000$dump_out$046;
  assign snapshot_packers$000$pack_in_$047 = snapshots$000$dump_out$047;
  assign snapshot_packers$000$pack_in_$048 = snapshots$000$dump_out$048;
  assign snapshot_packers$000$pack_in_$049 = snapshots$000$dump_out$049;
  assign snapshot_packers$000$pack_in_$050 = snapshots$000$dump_out$050;
  assign snapshot_packers$000$pack_in_$051 = snapshots$000$dump_out$051;
  assign snapshot_packers$000$pack_in_$052 = snapshots$000$dump_out$052;
  assign snapshot_packers$000$pack_in_$053 = snapshots$000$dump_out$053;
  assign snapshot_packers$000$pack_in_$054 = snapshots$000$dump_out$054;
  assign snapshot_packers$000$pack_in_$055 = snapshots$000$dump_out$055;
  assign snapshot_packers$000$pack_in_$056 = snapshots$000$dump_out$056;
  assign snapshot_packers$000$pack_in_$057 = snapshots$000$dump_out$057;
  assign snapshot_packers$000$pack_in_$058 = snapshots$000$dump_out$058;
  assign snapshot_packers$000$pack_in_$059 = snapshots$000$dump_out$059;
  assign snapshot_packers$000$pack_in_$060 = snapshots$000$dump_out$060;
  assign snapshot_packers$000$pack_in_$061 = snapshots$000$dump_out$061;
  assign snapshot_packers$000$pack_in_$062 = snapshots$000$dump_out$062;
  assign snapshot_packers$000$reset        = reset;
  assign snapshot_packers$001$clk          = clk;
  assign snapshot_packers$001$pack_in_$000 = snapshots$001$dump_out$000;
  assign snapshot_packers$001$pack_in_$001 = snapshots$001$dump_out$001;
  assign snapshot_packers$001$pack_in_$002 = snapshots$001$dump_out$002;
  assign snapshot_packers$001$pack_in_$003 = snapshots$001$dump_out$003;
  assign snapshot_packers$001$pack_in_$004 = snapshots$001$dump_out$004;
  assign snapshot_packers$001$pack_in_$005 = snapshots$001$dump_out$005;
  assign snapshot_packers$001$pack_in_$006 = snapshots$001$dump_out$006;
  assign snapshot_packers$001$pack_in_$007 = snapshots$001$dump_out$007;
  assign snapshot_packers$001$pack_in_$008 = snapshots$001$dump_out$008;
  assign snapshot_packers$001$pack_in_$009 = snapshots$001$dump_out$009;
  assign snapshot_packers$001$pack_in_$010 = snapshots$001$dump_out$010;
  assign snapshot_packers$001$pack_in_$011 = snapshots$001$dump_out$011;
  assign snapshot_packers$001$pack_in_$012 = snapshots$001$dump_out$012;
  assign snapshot_packers$001$pack_in_$013 = snapshots$001$dump_out$013;
  assign snapshot_packers$001$pack_in_$014 = snapshots$001$dump_out$014;
  assign snapshot_packers$001$pack_in_$015 = snapshots$001$dump_out$015;
  assign snapshot_packers$001$pack_in_$016 = snapshots$001$dump_out$016;
  assign snapshot_packers$001$pack_in_$017 = snapshots$001$dump_out$017;
  assign snapshot_packers$001$pack_in_$018 = snapshots$001$dump_out$018;
  assign snapshot_packers$001$pack_in_$019 = snapshots$001$dump_out$019;
  assign snapshot_packers$001$pack_in_$020 = snapshots$001$dump_out$020;
  assign snapshot_packers$001$pack_in_$021 = snapshots$001$dump_out$021;
  assign snapshot_packers$001$pack_in_$022 = snapshots$001$dump_out$022;
  assign snapshot_packers$001$pack_in_$023 = snapshots$001$dump_out$023;
  assign snapshot_packers$001$pack_in_$024 = snapshots$001$dump_out$024;
  assign snapshot_packers$001$pack_in_$025 = snapshots$001$dump_out$025;
  assign snapshot_packers$001$pack_in_$026 = snapshots$001$dump_out$026;
  assign snapshot_packers$001$pack_in_$027 = snapshots$001$dump_out$027;
  assign snapshot_packers$001$pack_in_$028 = snapshots$001$dump_out$028;
  assign snapshot_packers$001$pack_in_$029 = snapshots$001$dump_out$029;
  assign snapshot_packers$001$pack_in_$030 = snapshots$001$dump_out$030;
  assign snapshot_packers$001$pack_in_$031 = snapshots$001$dump_out$031;
  assign snapshot_packers$001$pack_in_$032 = snapshots$001$dump_out$032;
  assign snapshot_packers$001$pack_in_$033 = snapshots$001$dump_out$033;
  assign snapshot_packers$001$pack_in_$034 = snapshots$001$dump_out$034;
  assign snapshot_packers$001$pack_in_$035 = snapshots$001$dump_out$035;
  assign snapshot_packers$001$pack_in_$036 = snapshots$001$dump_out$036;
  assign snapshot_packers$001$pack_in_$037 = snapshots$001$dump_out$037;
  assign snapshot_packers$001$pack_in_$038 = snapshots$001$dump_out$038;
  assign snapshot_packers$001$pack_in_$039 = snapshots$001$dump_out$039;
  assign snapshot_packers$001$pack_in_$040 = snapshots$001$dump_out$040;
  assign snapshot_packers$001$pack_in_$041 = snapshots$001$dump_out$041;
  assign snapshot_packers$001$pack_in_$042 = snapshots$001$dump_out$042;
  assign snapshot_packers$001$pack_in_$043 = snapshots$001$dump_out$043;
  assign snapshot_packers$001$pack_in_$044 = snapshots$001$dump_out$044;
  assign snapshot_packers$001$pack_in_$045 = snapshots$001$dump_out$045;
  assign snapshot_packers$001$pack_in_$046 = snapshots$001$dump_out$046;
  assign snapshot_packers$001$pack_in_$047 = snapshots$001$dump_out$047;
  assign snapshot_packers$001$pack_in_$048 = snapshots$001$dump_out$048;
  assign snapshot_packers$001$pack_in_$049 = snapshots$001$dump_out$049;
  assign snapshot_packers$001$pack_in_$050 = snapshots$001$dump_out$050;
  assign snapshot_packers$001$pack_in_$051 = snapshots$001$dump_out$051;
  assign snapshot_packers$001$pack_in_$052 = snapshots$001$dump_out$052;
  assign snapshot_packers$001$pack_in_$053 = snapshots$001$dump_out$053;
  assign snapshot_packers$001$pack_in_$054 = snapshots$001$dump_out$054;
  assign snapshot_packers$001$pack_in_$055 = snapshots$001$dump_out$055;
  assign snapshot_packers$001$pack_in_$056 = snapshots$001$dump_out$056;
  assign snapshot_packers$001$pack_in_$057 = snapshots$001$dump_out$057;
  assign snapshot_packers$001$pack_in_$058 = snapshots$001$dump_out$058;
  assign snapshot_packers$001$pack_in_$059 = snapshots$001$dump_out$059;
  assign snapshot_packers$001$pack_in_$060 = snapshots$001$dump_out$060;
  assign snapshot_packers$001$pack_in_$061 = snapshots$001$dump_out$061;
  assign snapshot_packers$001$pack_in_$062 = snapshots$001$dump_out$062;
  assign snapshot_packers$001$reset        = reset;
  assign snapshots$000$clk                 = clk;
  assign snapshots$000$reset               = reset;
  assign snapshots$000$set_in_$000         = 1'd0;
  assign snapshots$000$set_in_$001         = 1'd0;
  assign snapshots$000$set_in_$002         = 1'd0;
  assign snapshots$000$set_in_$003         = 1'd0;
  assign snapshots$000$set_in_$004         = 1'd0;
  assign snapshots$000$set_in_$005         = 1'd0;
  assign snapshots$000$set_in_$006         = 1'd0;
  assign snapshots$000$set_in_$007         = 1'd0;
  assign snapshots$000$set_in_$008         = 1'd0;
  assign snapshots$000$set_in_$009         = 1'd0;
  assign snapshots$000$set_in_$010         = 1'd0;
  assign snapshots$000$set_in_$011         = 1'd0;
  assign snapshots$000$set_in_$012         = 1'd0;
  assign snapshots$000$set_in_$013         = 1'd0;
  assign snapshots$000$set_in_$014         = 1'd0;
  assign snapshots$000$set_in_$015         = 1'd0;
  assign snapshots$000$set_in_$016         = 1'd0;
  assign snapshots$000$set_in_$017         = 1'd0;
  assign snapshots$000$set_in_$018         = 1'd0;
  assign snapshots$000$set_in_$019         = 1'd0;
  assign snapshots$000$set_in_$020         = 1'd0;
  assign snapshots$000$set_in_$021         = 1'd0;
  assign snapshots$000$set_in_$022         = 1'd0;
  assign snapshots$000$set_in_$023         = 1'd0;
  assign snapshots$000$set_in_$024         = 1'd0;
  assign snapshots$000$set_in_$025         = 1'd0;
  assign snapshots$000$set_in_$026         = 1'd0;
  assign snapshots$000$set_in_$027         = 1'd0;
  assign snapshots$000$set_in_$028         = 1'd0;
  assign snapshots$000$set_in_$029         = 1'd0;
  assign snapshots$000$set_in_$030         = 1'd0;
  assign snapshots$000$set_in_$031         = 1'd0;
  assign snapshots$000$set_in_$032         = 1'd0;
  assign snapshots$000$set_in_$033         = 1'd0;
  assign snapshots$000$set_in_$034         = 1'd0;
  assign snapshots$000$set_in_$035         = 1'd0;
  assign snapshots$000$set_in_$036         = 1'd0;
  assign snapshots$000$set_in_$037         = 1'd0;
  assign snapshots$000$set_in_$038         = 1'd0;
  assign snapshots$000$set_in_$039         = 1'd0;
  assign snapshots$000$set_in_$040         = 1'd0;
  assign snapshots$000$set_in_$041         = 1'd0;
  assign snapshots$000$set_in_$042         = 1'd0;
  assign snapshots$000$set_in_$043         = 1'd0;
  assign snapshots$000$set_in_$044         = 1'd0;
  assign snapshots$000$set_in_$045         = 1'd0;
  assign snapshots$000$set_in_$046         = 1'd0;
  assign snapshots$000$set_in_$047         = 1'd0;
  assign snapshots$000$set_in_$048         = 1'd0;
  assign snapshots$000$set_in_$049         = 1'd0;
  assign snapshots$000$set_in_$050         = 1'd0;
  assign snapshots$000$set_in_$051         = 1'd0;
  assign snapshots$000$set_in_$052         = 1'd0;
  assign snapshots$000$set_in_$053         = 1'd0;
  assign snapshots$000$set_in_$054         = 1'd0;
  assign snapshots$000$set_in_$055         = 1'd0;
  assign snapshots$000$set_in_$056         = 1'd0;
  assign snapshots$000$set_in_$057         = 1'd0;
  assign snapshots$000$set_in_$058         = 1'd0;
  assign snapshots$000$set_in_$059         = 1'd0;
  assign snapshots$000$set_in_$060         = 1'd0;
  assign snapshots$000$set_in_$061         = 1'd0;
  assign snapshots$000$set_in_$062         = 1'd0;
  assign snapshots$000$write_addr$000      = alloc_index$000;
  assign snapshots$000$write_call$000      = alloc_call$000;
  assign snapshots$000$write_data$000      = 1'd1;
  assign snapshots$001$clk                 = clk;
  assign snapshots$001$reset               = reset;
  assign snapshots$001$set_in_$000         = 1'd0;
  assign snapshots$001$set_in_$001         = 1'd0;
  assign snapshots$001$set_in_$002         = 1'd0;
  assign snapshots$001$set_in_$003         = 1'd0;
  assign snapshots$001$set_in_$004         = 1'd0;
  assign snapshots$001$set_in_$005         = 1'd0;
  assign snapshots$001$set_in_$006         = 1'd0;
  assign snapshots$001$set_in_$007         = 1'd0;
  assign snapshots$001$set_in_$008         = 1'd0;
  assign snapshots$001$set_in_$009         = 1'd0;
  assign snapshots$001$set_in_$010         = 1'd0;
  assign snapshots$001$set_in_$011         = 1'd0;
  assign snapshots$001$set_in_$012         = 1'd0;
  assign snapshots$001$set_in_$013         = 1'd0;
  assign snapshots$001$set_in_$014         = 1'd0;
  assign snapshots$001$set_in_$015         = 1'd0;
  assign snapshots$001$set_in_$016         = 1'd0;
  assign snapshots$001$set_in_$017         = 1'd0;
  assign snapshots$001$set_in_$018         = 1'd0;
  assign snapshots$001$set_in_$019         = 1'd0;
  assign snapshots$001$set_in_$020         = 1'd0;
  assign snapshots$001$set_in_$021         = 1'd0;
  assign snapshots$001$set_in_$022         = 1'd0;
  assign snapshots$001$set_in_$023         = 1'd0;
  assign snapshots$001$set_in_$024         = 1'd0;
  assign snapshots$001$set_in_$025         = 1'd0;
  assign snapshots$001$set_in_$026         = 1'd0;
  assign snapshots$001$set_in_$027         = 1'd0;
  assign snapshots$001$set_in_$028         = 1'd0;
  assign snapshots$001$set_in_$029         = 1'd0;
  assign snapshots$001$set_in_$030         = 1'd0;
  assign snapshots$001$set_in_$031         = 1'd0;
  assign snapshots$001$set_in_$032         = 1'd0;
  assign snapshots$001$set_in_$033         = 1'd0;
  assign snapshots$001$set_in_$034         = 1'd0;
  assign snapshots$001$set_in_$035         = 1'd0;
  assign snapshots$001$set_in_$036         = 1'd0;
  assign snapshots$001$set_in_$037         = 1'd0;
  assign snapshots$001$set_in_$038         = 1'd0;
  assign snapshots$001$set_in_$039         = 1'd0;
  assign snapshots$001$set_in_$040         = 1'd0;
  assign snapshots$001$set_in_$041         = 1'd0;
  assign snapshots$001$set_in_$042         = 1'd0;
  assign snapshots$001$set_in_$043         = 1'd0;
  assign snapshots$001$set_in_$044         = 1'd0;
  assign snapshots$001$set_in_$045         = 1'd0;
  assign snapshots$001$set_in_$046         = 1'd0;
  assign snapshots$001$set_in_$047         = 1'd0;
  assign snapshots$001$set_in_$048         = 1'd0;
  assign snapshots$001$set_in_$049         = 1'd0;
  assign snapshots$001$set_in_$050         = 1'd0;
  assign snapshots$001$set_in_$051         = 1'd0;
  assign snapshots$001$set_in_$052         = 1'd0;
  assign snapshots$001$set_in_$053         = 1'd0;
  assign snapshots$001$set_in_$054         = 1'd0;
  assign snapshots$001$set_in_$055         = 1'd0;
  assign snapshots$001$set_in_$056         = 1'd0;
  assign snapshots$001$set_in_$057         = 1'd0;
  assign snapshots$001$set_in_$058         = 1'd0;
  assign snapshots$001$set_in_$059         = 1'd0;
  assign snapshots$001$set_in_$060         = 1'd0;
  assign snapshots$001$set_in_$061         = 1'd0;
  assign snapshots$001$set_in_$062         = 1'd0;
  assign snapshots$001$write_addr$000      = alloc_index$000;
  assign snapshots$001$write_call$000      = alloc_call$000;
  assign snapshots$001$write_data$000      = 1'd1;

  // array declarations
  logic    [   0:0] snapshots$set_call[0:1];
  assign snapshots$000$set_call = snapshots$set_call[  0];
  assign snapshots$001$set_call = snapshots$set_call[  1];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_reset_alloc_tracking_set_call(i=i):
  //         if s.reset_alloc_tracking_call and s.reset_alloc_tracking_target_id == i:
  //           s.snapshots[i].set_call.v = 1
  //         else:
  //           s.snapshots[i].set_call.v = 0

  // logic for handle_reset_alloc_tracking_set_call()
  always @ (*) begin
    if ((reset_alloc_tracking_call&&(reset_alloc_tracking_target_id == 0))) begin
      snapshots$set_call[0] = 1;
    end
    else begin
      snapshots$set_call[0] = 0;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_reset_alloc_tracking_set_call(i=i):
  //         if s.reset_alloc_tracking_call and s.reset_alloc_tracking_target_id == i:
  //           s.snapshots[i].set_call.v = 1
  //         else:
  //           s.snapshots[i].set_call.v = 0

  // logic for handle_reset_alloc_tracking_set_call()
  always @ (*) begin
    if ((reset_alloc_tracking_call&&(reset_alloc_tracking_target_id == 1))) begin
      snapshots$set_call[1] = 1;
    end
    else begin
      snapshots$set_call[1] = 0;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_revert_alloc():
  //       if s.reset_alloc_tracking_call and s.revert_allocs_call and s.reset_alloc_tracking_target_id == s.revert_allocs_source_id:
  //         s.free_list.release_call.v = 0
  //       else:
  //         s.free_list.release_call.v = s.revert_allocs_call

  // logic for handle_revert_alloc()
  always @ (*) begin
    if ((reset_alloc_tracking_call&&revert_allocs_call&&(reset_alloc_tracking_target_id == revert_allocs_source_id))) begin
      free_list$release_call = 0;
    end
    else begin
      free_list$release_call = revert_allocs_call;
    end
  end


endmodule // SnapshottingFreeList_0x68f914e32e2c4f6d

//-----------------------------------------------------------------------------
// RegisterFile_0x764ec1b6bf9dc34b
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.registerfile {"dtype": 1, "nregs": 63, "num_read_ports": 0, "num_write_ports": 1, "reset_values": null, "write_dump_bypass": true, "write_read_bypass": false}
// PyMTL: verilator_xinit = zeros
module RegisterFile_0x764ec1b6bf9dc34b
(
  input  logic [   0:0] clk,
  output logic [   0:0] dump_out$000,
  output logic [   0:0] dump_out$010,
  output logic [   0:0] dump_out$011,
  output logic [   0:0] dump_out$012,
  output logic [   0:0] dump_out$013,
  output logic [   0:0] dump_out$014,
  output logic [   0:0] dump_out$015,
  output logic [   0:0] dump_out$016,
  output logic [   0:0] dump_out$017,
  output logic [   0:0] dump_out$018,
  output logic [   0:0] dump_out$019,
  output logic [   0:0] dump_out$001,
  output logic [   0:0] dump_out$020,
  output logic [   0:0] dump_out$021,
  output logic [   0:0] dump_out$022,
  output logic [   0:0] dump_out$023,
  output logic [   0:0] dump_out$024,
  output logic [   0:0] dump_out$025,
  output logic [   0:0] dump_out$026,
  output logic [   0:0] dump_out$027,
  output logic [   0:0] dump_out$028,
  output logic [   0:0] dump_out$029,
  output logic [   0:0] dump_out$002,
  output logic [   0:0] dump_out$030,
  output logic [   0:0] dump_out$031,
  output logic [   0:0] dump_out$032,
  output logic [   0:0] dump_out$033,
  output logic [   0:0] dump_out$034,
  output logic [   0:0] dump_out$035,
  output logic [   0:0] dump_out$036,
  output logic [   0:0] dump_out$037,
  output logic [   0:0] dump_out$038,
  output logic [   0:0] dump_out$039,
  output logic [   0:0] dump_out$003,
  output logic [   0:0] dump_out$040,
  output logic [   0:0] dump_out$041,
  output logic [   0:0] dump_out$042,
  output logic [   0:0] dump_out$043,
  output logic [   0:0] dump_out$044,
  output logic [   0:0] dump_out$045,
  output logic [   0:0] dump_out$046,
  output logic [   0:0] dump_out$047,
  output logic [   0:0] dump_out$048,
  output logic [   0:0] dump_out$049,
  output logic [   0:0] dump_out$004,
  output logic [   0:0] dump_out$050,
  output logic [   0:0] dump_out$051,
  output logic [   0:0] dump_out$052,
  output logic [   0:0] dump_out$053,
  output logic [   0:0] dump_out$054,
  output logic [   0:0] dump_out$055,
  output logic [   0:0] dump_out$056,
  output logic [   0:0] dump_out$057,
  output logic [   0:0] dump_out$058,
  output logic [   0:0] dump_out$059,
  output logic [   0:0] dump_out$005,
  output logic [   0:0] dump_out$060,
  output logic [   0:0] dump_out$061,
  output logic [   0:0] dump_out$062,
  output logic [   0:0] dump_out$006,
  output logic [   0:0] dump_out$007,
  output logic [   0:0] dump_out$008,
  output logic [   0:0] dump_out$009,
  input  logic [   0:0] reset,
  input  logic [   0:0] set_call,
  input  logic [   0:0] set_in_$000,
  input  logic [   0:0] set_in_$010,
  input  logic [   0:0] set_in_$011,
  input  logic [   0:0] set_in_$012,
  input  logic [   0:0] set_in_$013,
  input  logic [   0:0] set_in_$014,
  input  logic [   0:0] set_in_$015,
  input  logic [   0:0] set_in_$016,
  input  logic [   0:0] set_in_$017,
  input  logic [   0:0] set_in_$018,
  input  logic [   0:0] set_in_$019,
  input  logic [   0:0] set_in_$001,
  input  logic [   0:0] set_in_$020,
  input  logic [   0:0] set_in_$021,
  input  logic [   0:0] set_in_$022,
  input  logic [   0:0] set_in_$023,
  input  logic [   0:0] set_in_$024,
  input  logic [   0:0] set_in_$025,
  input  logic [   0:0] set_in_$026,
  input  logic [   0:0] set_in_$027,
  input  logic [   0:0] set_in_$028,
  input  logic [   0:0] set_in_$029,
  input  logic [   0:0] set_in_$002,
  input  logic [   0:0] set_in_$030,
  input  logic [   0:0] set_in_$031,
  input  logic [   0:0] set_in_$032,
  input  logic [   0:0] set_in_$033,
  input  logic [   0:0] set_in_$034,
  input  logic [   0:0] set_in_$035,
  input  logic [   0:0] set_in_$036,
  input  logic [   0:0] set_in_$037,
  input  logic [   0:0] set_in_$038,
  input  logic [   0:0] set_in_$039,
  input  logic [   0:0] set_in_$003,
  input  logic [   0:0] set_in_$040,
  input  logic [   0:0] set_in_$041,
  input  logic [   0:0] set_in_$042,
  input  logic [   0:0] set_in_$043,
  input  logic [   0:0] set_in_$044,
  input  logic [   0:0] set_in_$045,
  input  logic [   0:0] set_in_$046,
  input  logic [   0:0] set_in_$047,
  input  logic [   0:0] set_in_$048,
  input  logic [   0:0] set_in_$049,
  input  logic [   0:0] set_in_$004,
  input  logic [   0:0] set_in_$050,
  input  logic [   0:0] set_in_$051,
  input  logic [   0:0] set_in_$052,
  input  logic [   0:0] set_in_$053,
  input  logic [   0:0] set_in_$054,
  input  logic [   0:0] set_in_$055,
  input  logic [   0:0] set_in_$056,
  input  logic [   0:0] set_in_$057,
  input  logic [   0:0] set_in_$058,
  input  logic [   0:0] set_in_$059,
  input  logic [   0:0] set_in_$005,
  input  logic [   0:0] set_in_$060,
  input  logic [   0:0] set_in_$061,
  input  logic [   0:0] set_in_$062,
  input  logic [   0:0] set_in_$006,
  input  logic [   0:0] set_in_$007,
  input  logic [   0:0] set_in_$008,
  input  logic [   0:0] set_in_$009,
  input  logic [   5:0] write_addr$000,
  input  logic [   0:0] write_call$000,
  input  logic [   0:0] write_data$000
);

  // logic declarations
  logic   [   0:0] write_inc$000;
  logic   [   0:0] write_inc$001;
  logic   [   0:0] write_inc$002;
  logic   [   0:0] write_inc$003;
  logic   [   0:0] write_inc$004;
  logic   [   0:0] write_inc$005;
  logic   [   0:0] write_inc$006;
  logic   [   0:0] write_inc$007;
  logic   [   0:0] write_inc$008;
  logic   [   0:0] write_inc$009;
  logic   [   0:0] write_inc$010;
  logic   [   0:0] write_inc$011;
  logic   [   0:0] write_inc$012;
  logic   [   0:0] write_inc$013;
  logic   [   0:0] write_inc$014;
  logic   [   0:0] write_inc$015;
  logic   [   0:0] write_inc$016;
  logic   [   0:0] write_inc$017;
  logic   [   0:0] write_inc$018;
  logic   [   0:0] write_inc$019;
  logic   [   0:0] write_inc$020;
  logic   [   0:0] write_inc$021;
  logic   [   0:0] write_inc$022;
  logic   [   0:0] write_inc$023;
  logic   [   0:0] write_inc$024;
  logic   [   0:0] write_inc$025;
  logic   [   0:0] write_inc$026;
  logic   [   0:0] write_inc$027;
  logic   [   0:0] write_inc$028;
  logic   [   0:0] write_inc$029;
  logic   [   0:0] write_inc$030;
  logic   [   0:0] write_inc$031;
  logic   [   0:0] write_inc$032;
  logic   [   0:0] write_inc$033;
  logic   [   0:0] write_inc$034;
  logic   [   0:0] write_inc$035;
  logic   [   0:0] write_inc$036;
  logic   [   0:0] write_inc$037;
  logic   [   0:0] write_inc$038;
  logic   [   0:0] write_inc$039;
  logic   [   0:0] write_inc$040;
  logic   [   0:0] write_inc$041;
  logic   [   0:0] write_inc$042;
  logic   [   0:0] write_inc$043;
  logic   [   0:0] write_inc$044;
  logic   [   0:0] write_inc$045;
  logic   [   0:0] write_inc$046;
  logic   [   0:0] write_inc$047;
  logic   [   0:0] write_inc$048;
  logic   [   0:0] write_inc$049;
  logic   [   0:0] write_inc$050;
  logic   [   0:0] write_inc$051;
  logic   [   0:0] write_inc$052;
  logic   [   0:0] write_inc$053;
  logic   [   0:0] write_inc$054;
  logic   [   0:0] write_inc$055;
  logic   [   0:0] write_inc$056;
  logic   [   0:0] write_inc$057;
  logic   [   0:0] write_inc$058;
  logic   [   0:0] write_inc$059;
  logic   [   0:0] write_inc$060;
  logic   [   0:0] write_inc$061;
  logic   [   0:0] write_inc$062;
  logic   [   0:0] after_set$000;
  logic   [   0:0] after_set$001;
  logic   [   0:0] after_set$002;
  logic   [   0:0] after_set$003;
  logic   [   0:0] after_set$004;
  logic   [   0:0] after_set$005;
  logic   [   0:0] after_set$006;
  logic   [   0:0] after_set$007;
  logic   [   0:0] after_set$008;
  logic   [   0:0] after_set$009;
  logic   [   0:0] after_set$010;
  logic   [   0:0] after_set$011;
  logic   [   0:0] after_set$012;
  logic   [   0:0] after_set$013;
  logic   [   0:0] after_set$014;
  logic   [   0:0] after_set$015;
  logic   [   0:0] after_set$016;
  logic   [   0:0] after_set$017;
  logic   [   0:0] after_set$018;
  logic   [   0:0] after_set$019;
  logic   [   0:0] after_set$020;
  logic   [   0:0] after_set$021;
  logic   [   0:0] after_set$022;
  logic   [   0:0] after_set$023;
  logic   [   0:0] after_set$024;
  logic   [   0:0] after_set$025;
  logic   [   0:0] after_set$026;
  logic   [   0:0] after_set$027;
  logic   [   0:0] after_set$028;
  logic   [   0:0] after_set$029;
  logic   [   0:0] after_set$030;
  logic   [   0:0] after_set$031;
  logic   [   0:0] after_set$032;
  logic   [   0:0] after_set$033;
  logic   [   0:0] after_set$034;
  logic   [   0:0] after_set$035;
  logic   [   0:0] after_set$036;
  logic   [   0:0] after_set$037;
  logic   [   0:0] after_set$038;
  logic   [   0:0] after_set$039;
  logic   [   0:0] after_set$040;
  logic   [   0:0] after_set$041;
  logic   [   0:0] after_set$042;
  logic   [   0:0] after_set$043;
  logic   [   0:0] after_set$044;
  logic   [   0:0] after_set$045;
  logic   [   0:0] after_set$046;
  logic   [   0:0] after_set$047;
  logic   [   0:0] after_set$048;
  logic   [   0:0] after_set$049;
  logic   [   0:0] after_set$050;
  logic   [   0:0] after_set$051;
  logic   [   0:0] after_set$052;
  logic   [   0:0] after_set$053;
  logic   [   0:0] after_set$054;
  logic   [   0:0] after_set$055;
  logic   [   0:0] after_set$056;
  logic   [   0:0] after_set$057;
  logic   [   0:0] after_set$058;
  logic   [   0:0] after_set$059;
  logic   [   0:0] after_set$060;
  logic   [   0:0] after_set$061;
  logic   [   0:0] after_set$062;
  logic   [   0:0] regs$000;
  logic   [   0:0] regs$001;
  logic   [   0:0] regs$002;
  logic   [   0:0] regs$003;
  logic   [   0:0] regs$004;
  logic   [   0:0] regs$005;
  logic   [   0:0] regs$006;
  logic   [   0:0] regs$007;
  logic   [   0:0] regs$008;
  logic   [   0:0] regs$009;
  logic   [   0:0] regs$010;
  logic   [   0:0] regs$011;
  logic   [   0:0] regs$012;
  logic   [   0:0] regs$013;
  logic   [   0:0] regs$014;
  logic   [   0:0] regs$015;
  logic   [   0:0] regs$016;
  logic   [   0:0] regs$017;
  logic   [   0:0] regs$018;
  logic   [   0:0] regs$019;
  logic   [   0:0] regs$020;
  logic   [   0:0] regs$021;
  logic   [   0:0] regs$022;
  logic   [   0:0] regs$023;
  logic   [   0:0] regs$024;
  logic   [   0:0] regs$025;
  logic   [   0:0] regs$026;
  logic   [   0:0] regs$027;
  logic   [   0:0] regs$028;
  logic   [   0:0] regs$029;
  logic   [   0:0] regs$030;
  logic   [   0:0] regs$031;
  logic   [   0:0] regs$032;
  logic   [   0:0] regs$033;
  logic   [   0:0] regs$034;
  logic   [   0:0] regs$035;
  logic   [   0:0] regs$036;
  logic   [   0:0] regs$037;
  logic   [   0:0] regs$038;
  logic   [   0:0] regs$039;
  logic   [   0:0] regs$040;
  logic   [   0:0] regs$041;
  logic   [   0:0] regs$042;
  logic   [   0:0] regs$043;
  logic   [   0:0] regs$044;
  logic   [   0:0] regs$045;
  logic   [   0:0] regs$046;
  logic   [   0:0] regs$047;
  logic   [   0:0] regs$048;
  logic   [   0:0] regs$049;
  logic   [   0:0] regs$050;
  logic   [   0:0] regs$051;
  logic   [   0:0] regs$052;
  logic   [   0:0] regs$053;
  logic   [   0:0] regs$054;
  logic   [   0:0] regs$055;
  logic   [   0:0] regs$056;
  logic   [   0:0] regs$057;
  logic   [   0:0] regs$058;
  logic   [   0:0] regs$059;
  logic   [   0:0] regs$060;
  logic   [   0:0] regs$061;
  logic   [   0:0] regs$062;
  logic   [   0:0] after_write$000;
  logic   [   0:0] after_write$001;
  logic   [   0:0] after_write$002;
  logic   [   0:0] after_write$003;
  logic   [   0:0] after_write$004;
  logic   [   0:0] after_write$005;
  logic   [   0:0] after_write$006;
  logic   [   0:0] after_write$007;
  logic   [   0:0] after_write$008;
  logic   [   0:0] after_write$009;
  logic   [   0:0] after_write$010;
  logic   [   0:0] after_write$011;
  logic   [   0:0] after_write$012;
  logic   [   0:0] after_write$013;
  logic   [   0:0] after_write$014;
  logic   [   0:0] after_write$015;
  logic   [   0:0] after_write$016;
  logic   [   0:0] after_write$017;
  logic   [   0:0] after_write$018;
  logic   [   0:0] after_write$019;
  logic   [   0:0] after_write$020;
  logic   [   0:0] after_write$021;
  logic   [   0:0] after_write$022;
  logic   [   0:0] after_write$023;
  logic   [   0:0] after_write$024;
  logic   [   0:0] after_write$025;
  logic   [   0:0] after_write$026;
  logic   [   0:0] after_write$027;
  logic   [   0:0] after_write$028;
  logic   [   0:0] after_write$029;
  logic   [   0:0] after_write$030;
  logic   [   0:0] after_write$031;
  logic   [   0:0] after_write$032;
  logic   [   0:0] after_write$033;
  logic   [   0:0] after_write$034;
  logic   [   0:0] after_write$035;
  logic   [   0:0] after_write$036;
  logic   [   0:0] after_write$037;
  logic   [   0:0] after_write$038;
  logic   [   0:0] after_write$039;
  logic   [   0:0] after_write$040;
  logic   [   0:0] after_write$041;
  logic   [   0:0] after_write$042;
  logic   [   0:0] after_write$043;
  logic   [   0:0] after_write$044;
  logic   [   0:0] after_write$045;
  logic   [   0:0] after_write$046;
  logic   [   0:0] after_write$047;
  logic   [   0:0] after_write$048;
  logic   [   0:0] after_write$049;
  logic   [   0:0] after_write$050;
  logic   [   0:0] after_write$051;
  logic   [   0:0] after_write$052;
  logic   [   0:0] after_write$053;
  logic   [   0:0] after_write$054;
  logic   [   0:0] after_write$055;
  logic   [   0:0] after_write$056;
  logic   [   0:0] after_write$057;
  logic   [   0:0] after_write$058;
  logic   [   0:0] after_write$059;
  logic   [   0:0] after_write$060;
  logic   [   0:0] after_write$061;
  logic   [   0:0] after_write$062;


  // signal connections
  assign dump_out$000 = after_write$000;
  assign dump_out$001 = after_write$001;
  assign dump_out$002 = after_write$002;
  assign dump_out$003 = after_write$003;
  assign dump_out$004 = after_write$004;
  assign dump_out$005 = after_write$005;
  assign dump_out$006 = after_write$006;
  assign dump_out$007 = after_write$007;
  assign dump_out$008 = after_write$008;
  assign dump_out$009 = after_write$009;
  assign dump_out$010 = after_write$010;
  assign dump_out$011 = after_write$011;
  assign dump_out$012 = after_write$012;
  assign dump_out$013 = after_write$013;
  assign dump_out$014 = after_write$014;
  assign dump_out$015 = after_write$015;
  assign dump_out$016 = after_write$016;
  assign dump_out$017 = after_write$017;
  assign dump_out$018 = after_write$018;
  assign dump_out$019 = after_write$019;
  assign dump_out$020 = after_write$020;
  assign dump_out$021 = after_write$021;
  assign dump_out$022 = after_write$022;
  assign dump_out$023 = after_write$023;
  assign dump_out$024 = after_write$024;
  assign dump_out$025 = after_write$025;
  assign dump_out$026 = after_write$026;
  assign dump_out$027 = after_write$027;
  assign dump_out$028 = after_write$028;
  assign dump_out$029 = after_write$029;
  assign dump_out$030 = after_write$030;
  assign dump_out$031 = after_write$031;
  assign dump_out$032 = after_write$032;
  assign dump_out$033 = after_write$033;
  assign dump_out$034 = after_write$034;
  assign dump_out$035 = after_write$035;
  assign dump_out$036 = after_write$036;
  assign dump_out$037 = after_write$037;
  assign dump_out$038 = after_write$038;
  assign dump_out$039 = after_write$039;
  assign dump_out$040 = after_write$040;
  assign dump_out$041 = after_write$041;
  assign dump_out$042 = after_write$042;
  assign dump_out$043 = after_write$043;
  assign dump_out$044 = after_write$044;
  assign dump_out$045 = after_write$045;
  assign dump_out$046 = after_write$046;
  assign dump_out$047 = after_write$047;
  assign dump_out$048 = after_write$048;
  assign dump_out$049 = after_write$049;
  assign dump_out$050 = after_write$050;
  assign dump_out$051 = after_write$051;
  assign dump_out$052 = after_write$052;
  assign dump_out$053 = after_write$053;
  assign dump_out$054 = after_write$054;
  assign dump_out$055 = after_write$055;
  assign dump_out$056 = after_write$056;
  assign dump_out$057 = after_write$057;
  assign dump_out$058 = after_write$058;
  assign dump_out$059 = after_write$059;
  assign dump_out$060 = after_write$060;
  assign dump_out$061 = after_write$061;
  assign dump_out$062 = after_write$062;

  // array declarations
  logic    [   0:0] after_set[0:62];
  assign after_set$000 = after_set[  0];
  assign after_set$001 = after_set[  1];
  assign after_set$002 = after_set[  2];
  assign after_set$003 = after_set[  3];
  assign after_set$004 = after_set[  4];
  assign after_set$005 = after_set[  5];
  assign after_set$006 = after_set[  6];
  assign after_set$007 = after_set[  7];
  assign after_set$008 = after_set[  8];
  assign after_set$009 = after_set[  9];
  assign after_set$010 = after_set[ 10];
  assign after_set$011 = after_set[ 11];
  assign after_set$012 = after_set[ 12];
  assign after_set$013 = after_set[ 13];
  assign after_set$014 = after_set[ 14];
  assign after_set$015 = after_set[ 15];
  assign after_set$016 = after_set[ 16];
  assign after_set$017 = after_set[ 17];
  assign after_set$018 = after_set[ 18];
  assign after_set$019 = after_set[ 19];
  assign after_set$020 = after_set[ 20];
  assign after_set$021 = after_set[ 21];
  assign after_set$022 = after_set[ 22];
  assign after_set$023 = after_set[ 23];
  assign after_set$024 = after_set[ 24];
  assign after_set$025 = after_set[ 25];
  assign after_set$026 = after_set[ 26];
  assign after_set$027 = after_set[ 27];
  assign after_set$028 = after_set[ 28];
  assign after_set$029 = after_set[ 29];
  assign after_set$030 = after_set[ 30];
  assign after_set$031 = after_set[ 31];
  assign after_set$032 = after_set[ 32];
  assign after_set$033 = after_set[ 33];
  assign after_set$034 = after_set[ 34];
  assign after_set$035 = after_set[ 35];
  assign after_set$036 = after_set[ 36];
  assign after_set$037 = after_set[ 37];
  assign after_set$038 = after_set[ 38];
  assign after_set$039 = after_set[ 39];
  assign after_set$040 = after_set[ 40];
  assign after_set$041 = after_set[ 41];
  assign after_set$042 = after_set[ 42];
  assign after_set$043 = after_set[ 43];
  assign after_set$044 = after_set[ 44];
  assign after_set$045 = after_set[ 45];
  assign after_set$046 = after_set[ 46];
  assign after_set$047 = after_set[ 47];
  assign after_set$048 = after_set[ 48];
  assign after_set$049 = after_set[ 49];
  assign after_set$050 = after_set[ 50];
  assign after_set$051 = after_set[ 51];
  assign after_set$052 = after_set[ 52];
  assign after_set$053 = after_set[ 53];
  assign after_set$054 = after_set[ 54];
  assign after_set$055 = after_set[ 55];
  assign after_set$056 = after_set[ 56];
  assign after_set$057 = after_set[ 57];
  assign after_set$058 = after_set[ 58];
  assign after_set$059 = after_set[ 59];
  assign after_set$060 = after_set[ 60];
  assign after_set$061 = after_set[ 61];
  assign after_set$062 = after_set[ 62];
  logic    [   0:0] after_write[0:62];
  assign after_write$000 = after_write[  0];
  assign after_write$001 = after_write[  1];
  assign after_write$002 = after_write[  2];
  assign after_write$003 = after_write[  3];
  assign after_write$004 = after_write[  4];
  assign after_write$005 = after_write[  5];
  assign after_write$006 = after_write[  6];
  assign after_write$007 = after_write[  7];
  assign after_write$008 = after_write[  8];
  assign after_write$009 = after_write[  9];
  assign after_write$010 = after_write[ 10];
  assign after_write$011 = after_write[ 11];
  assign after_write$012 = after_write[ 12];
  assign after_write$013 = after_write[ 13];
  assign after_write$014 = after_write[ 14];
  assign after_write$015 = after_write[ 15];
  assign after_write$016 = after_write[ 16];
  assign after_write$017 = after_write[ 17];
  assign after_write$018 = after_write[ 18];
  assign after_write$019 = after_write[ 19];
  assign after_write$020 = after_write[ 20];
  assign after_write$021 = after_write[ 21];
  assign after_write$022 = after_write[ 22];
  assign after_write$023 = after_write[ 23];
  assign after_write$024 = after_write[ 24];
  assign after_write$025 = after_write[ 25];
  assign after_write$026 = after_write[ 26];
  assign after_write$027 = after_write[ 27];
  assign after_write$028 = after_write[ 28];
  assign after_write$029 = after_write[ 29];
  assign after_write$030 = after_write[ 30];
  assign after_write$031 = after_write[ 31];
  assign after_write$032 = after_write[ 32];
  assign after_write$033 = after_write[ 33];
  assign after_write$034 = after_write[ 34];
  assign after_write$035 = after_write[ 35];
  assign after_write$036 = after_write[ 36];
  assign after_write$037 = after_write[ 37];
  assign after_write$038 = after_write[ 38];
  assign after_write$039 = after_write[ 39];
  assign after_write$040 = after_write[ 40];
  assign after_write$041 = after_write[ 41];
  assign after_write$042 = after_write[ 42];
  assign after_write$043 = after_write[ 43];
  assign after_write$044 = after_write[ 44];
  assign after_write$045 = after_write[ 45];
  assign after_write$046 = after_write[ 46];
  assign after_write$047 = after_write[ 47];
  assign after_write$048 = after_write[ 48];
  assign after_write$049 = after_write[ 49];
  assign after_write$050 = after_write[ 50];
  assign after_write$051 = after_write[ 51];
  assign after_write$052 = after_write[ 52];
  assign after_write$053 = after_write[ 53];
  assign after_write$054 = after_write[ 54];
  assign after_write$055 = after_write[ 55];
  assign after_write$056 = after_write[ 56];
  assign after_write$057 = after_write[ 57];
  assign after_write$058 = after_write[ 58];
  assign after_write$059 = after_write[ 59];
  assign after_write$060 = after_write[ 60];
  assign after_write$061 = after_write[ 61];
  assign after_write$062 = after_write[ 62];
  logic    [   0:0] regs[0:62];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  assign regs$002 = regs[  2];
  assign regs$003 = regs[  3];
  assign regs$004 = regs[  4];
  assign regs$005 = regs[  5];
  assign regs$006 = regs[  6];
  assign regs$007 = regs[  7];
  assign regs$008 = regs[  8];
  assign regs$009 = regs[  9];
  assign regs$010 = regs[ 10];
  assign regs$011 = regs[ 11];
  assign regs$012 = regs[ 12];
  assign regs$013 = regs[ 13];
  assign regs$014 = regs[ 14];
  assign regs$015 = regs[ 15];
  assign regs$016 = regs[ 16];
  assign regs$017 = regs[ 17];
  assign regs$018 = regs[ 18];
  assign regs$019 = regs[ 19];
  assign regs$020 = regs[ 20];
  assign regs$021 = regs[ 21];
  assign regs$022 = regs[ 22];
  assign regs$023 = regs[ 23];
  assign regs$024 = regs[ 24];
  assign regs$025 = regs[ 25];
  assign regs$026 = regs[ 26];
  assign regs$027 = regs[ 27];
  assign regs$028 = regs[ 28];
  assign regs$029 = regs[ 29];
  assign regs$030 = regs[ 30];
  assign regs$031 = regs[ 31];
  assign regs$032 = regs[ 32];
  assign regs$033 = regs[ 33];
  assign regs$034 = regs[ 34];
  assign regs$035 = regs[ 35];
  assign regs$036 = regs[ 36];
  assign regs$037 = regs[ 37];
  assign regs$038 = regs[ 38];
  assign regs$039 = regs[ 39];
  assign regs$040 = regs[ 40];
  assign regs$041 = regs[ 41];
  assign regs$042 = regs[ 42];
  assign regs$043 = regs[ 43];
  assign regs$044 = regs[ 44];
  assign regs$045 = regs[ 45];
  assign regs$046 = regs[ 46];
  assign regs$047 = regs[ 47];
  assign regs$048 = regs[ 48];
  assign regs$049 = regs[ 49];
  assign regs$050 = regs[ 50];
  assign regs$051 = regs[ 51];
  assign regs$052 = regs[ 52];
  assign regs$053 = regs[ 53];
  assign regs$054 = regs[ 54];
  assign regs$055 = regs[ 55];
  assign regs$056 = regs[ 56];
  assign regs$057 = regs[ 57];
  assign regs$058 = regs[ 58];
  assign regs$059 = regs[ 59];
  assign regs$060 = regs[ 60];
  assign regs$061 = regs[ 61];
  assign regs$062 = regs[ 62];
  logic   [   0:0] set_in_[0:62];
  assign set_in_[  0] = set_in_$000;
  assign set_in_[  1] = set_in_$001;
  assign set_in_[  2] = set_in_$002;
  assign set_in_[  3] = set_in_$003;
  assign set_in_[  4] = set_in_$004;
  assign set_in_[  5] = set_in_$005;
  assign set_in_[  6] = set_in_$006;
  assign set_in_[  7] = set_in_$007;
  assign set_in_[  8] = set_in_$008;
  assign set_in_[  9] = set_in_$009;
  assign set_in_[ 10] = set_in_$010;
  assign set_in_[ 11] = set_in_$011;
  assign set_in_[ 12] = set_in_$012;
  assign set_in_[ 13] = set_in_$013;
  assign set_in_[ 14] = set_in_$014;
  assign set_in_[ 15] = set_in_$015;
  assign set_in_[ 16] = set_in_$016;
  assign set_in_[ 17] = set_in_$017;
  assign set_in_[ 18] = set_in_$018;
  assign set_in_[ 19] = set_in_$019;
  assign set_in_[ 20] = set_in_$020;
  assign set_in_[ 21] = set_in_$021;
  assign set_in_[ 22] = set_in_$022;
  assign set_in_[ 23] = set_in_$023;
  assign set_in_[ 24] = set_in_$024;
  assign set_in_[ 25] = set_in_$025;
  assign set_in_[ 26] = set_in_$026;
  assign set_in_[ 27] = set_in_$027;
  assign set_in_[ 28] = set_in_$028;
  assign set_in_[ 29] = set_in_$029;
  assign set_in_[ 30] = set_in_$030;
  assign set_in_[ 31] = set_in_$031;
  assign set_in_[ 32] = set_in_$032;
  assign set_in_[ 33] = set_in_$033;
  assign set_in_[ 34] = set_in_$034;
  assign set_in_[ 35] = set_in_$035;
  assign set_in_[ 36] = set_in_$036;
  assign set_in_[ 37] = set_in_$037;
  assign set_in_[ 38] = set_in_$038;
  assign set_in_[ 39] = set_in_$039;
  assign set_in_[ 40] = set_in_$040;
  assign set_in_[ 41] = set_in_$041;
  assign set_in_[ 42] = set_in_$042;
  assign set_in_[ 43] = set_in_$043;
  assign set_in_[ 44] = set_in_$044;
  assign set_in_[ 45] = set_in_$045;
  assign set_in_[ 46] = set_in_$046;
  assign set_in_[ 47] = set_in_$047;
  assign set_in_[ 48] = set_in_$048;
  assign set_in_[ 49] = set_in_$049;
  assign set_in_[ 50] = set_in_$050;
  assign set_in_[ 51] = set_in_$051;
  assign set_in_[ 52] = set_in_$052;
  assign set_in_[ 53] = set_in_$053;
  assign set_in_[ 54] = set_in_$054;
  assign set_in_[ 55] = set_in_$055;
  assign set_in_[ 56] = set_in_$056;
  assign set_in_[ 57] = set_in_$057;
  assign set_in_[ 58] = set_in_$058;
  assign set_in_[ 59] = set_in_$059;
  assign set_in_[ 60] = set_in_$060;
  assign set_in_[ 61] = set_in_$061;
  assign set_in_[ 62] = set_in_$062;
  logic   [   5:0] write_addr[0:0];
  assign write_addr[  0] = write_addr$000;
  logic   [   0:0] write_call[0:0];
  assign write_call[  0] = write_call$000;
  logic   [   0:0] write_data[0:0];
  assign write_data[  0] = write_data$000;
  logic    [   0:0] write_inc[0:62];
  assign write_inc$000 = write_inc[  0];
  assign write_inc$001 = write_inc[  1];
  assign write_inc$002 = write_inc[  2];
  assign write_inc$003 = write_inc[  3];
  assign write_inc$004 = write_inc[  4];
  assign write_inc$005 = write_inc[  5];
  assign write_inc$006 = write_inc[  6];
  assign write_inc$007 = write_inc[  7];
  assign write_inc$008 = write_inc[  8];
  assign write_inc$009 = write_inc[  9];
  assign write_inc$010 = write_inc[ 10];
  assign write_inc$011 = write_inc[ 11];
  assign write_inc$012 = write_inc[ 12];
  assign write_inc$013 = write_inc[ 13];
  assign write_inc$014 = write_inc[ 14];
  assign write_inc$015 = write_inc[ 15];
  assign write_inc$016 = write_inc[ 16];
  assign write_inc$017 = write_inc[ 17];
  assign write_inc$018 = write_inc[ 18];
  assign write_inc$019 = write_inc[ 19];
  assign write_inc$020 = write_inc[ 20];
  assign write_inc$021 = write_inc[ 21];
  assign write_inc$022 = write_inc[ 22];
  assign write_inc$023 = write_inc[ 23];
  assign write_inc$024 = write_inc[ 24];
  assign write_inc$025 = write_inc[ 25];
  assign write_inc$026 = write_inc[ 26];
  assign write_inc$027 = write_inc[ 27];
  assign write_inc$028 = write_inc[ 28];
  assign write_inc$029 = write_inc[ 29];
  assign write_inc$030 = write_inc[ 30];
  assign write_inc$031 = write_inc[ 31];
  assign write_inc$032 = write_inc[ 32];
  assign write_inc$033 = write_inc[ 33];
  assign write_inc$034 = write_inc[ 34];
  assign write_inc$035 = write_inc[ 35];
  assign write_inc$036 = write_inc[ 36];
  assign write_inc$037 = write_inc[ 37];
  assign write_inc$038 = write_inc[ 38];
  assign write_inc$039 = write_inc[ 39];
  assign write_inc$040 = write_inc[ 40];
  assign write_inc$041 = write_inc[ 41];
  assign write_inc$042 = write_inc[ 42];
  assign write_inc$043 = write_inc[ 43];
  assign write_inc$044 = write_inc[ 44];
  assign write_inc$045 = write_inc[ 45];
  assign write_inc$046 = write_inc[ 46];
  assign write_inc$047 = write_inc[ 47];
  assign write_inc$048 = write_inc[ 48];
  assign write_inc$049 = write_inc[ 49];
  assign write_inc$050 = write_inc[ 50];
  assign write_inc$051 = write_inc[ 51];
  assign write_inc$052 = write_inc[ 52];
  assign write_inc$053 = write_inc[ 53];
  assign write_inc$054 = write_inc[ 54];
  assign write_inc$055 = write_inc[ 55];
  assign write_inc$056 = write_inc[ 56];
  assign write_inc$057 = write_inc[ 57];
  assign write_inc$058 = write_inc[ 58];
  assign write_inc$059 = write_inc[ 59];
  assign write_inc$060 = write_inc[ 60];
  assign write_inc$061 = write_inc[ 61];
  assign write_inc$062 = write_inc[ 62];

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[0] <= 0;
    end
    else begin
      regs[0] <= after_set[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[1] <= 0;
    end
    else begin
      regs[1] <= after_set[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[2] <= 0;
    end
    else begin
      regs[2] <= after_set[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[3] <= 0;
    end
    else begin
      regs[3] <= after_set[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[4] <= 0;
    end
    else begin
      regs[4] <= after_set[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[5] <= 0;
    end
    else begin
      regs[5] <= after_set[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[6] <= 0;
    end
    else begin
      regs[6] <= after_set[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[7] <= 0;
    end
    else begin
      regs[7] <= after_set[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[8] <= 0;
    end
    else begin
      regs[8] <= after_set[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[9] <= 0;
    end
    else begin
      regs[9] <= after_set[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[10] <= 0;
    end
    else begin
      regs[10] <= after_set[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[11] <= 0;
    end
    else begin
      regs[11] <= after_set[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[12] <= 0;
    end
    else begin
      regs[12] <= after_set[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[13] <= 0;
    end
    else begin
      regs[13] <= after_set[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[14] <= 0;
    end
    else begin
      regs[14] <= after_set[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[15] <= 0;
    end
    else begin
      regs[15] <= after_set[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[16] <= 0;
    end
    else begin
      regs[16] <= after_set[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[17] <= 0;
    end
    else begin
      regs[17] <= after_set[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[18] <= 0;
    end
    else begin
      regs[18] <= after_set[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[19] <= 0;
    end
    else begin
      regs[19] <= after_set[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[20] <= 0;
    end
    else begin
      regs[20] <= after_set[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[21] <= 0;
    end
    else begin
      regs[21] <= after_set[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[22] <= 0;
    end
    else begin
      regs[22] <= after_set[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[23] <= 0;
    end
    else begin
      regs[23] <= after_set[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[24] <= 0;
    end
    else begin
      regs[24] <= after_set[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[25] <= 0;
    end
    else begin
      regs[25] <= after_set[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[26] <= 0;
    end
    else begin
      regs[26] <= after_set[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[27] <= 0;
    end
    else begin
      regs[27] <= after_set[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[28] <= 0;
    end
    else begin
      regs[28] <= after_set[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[29] <= 0;
    end
    else begin
      regs[29] <= after_set[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[30] <= 0;
    end
    else begin
      regs[30] <= after_set[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[31] <= 0;
    end
    else begin
      regs[31] <= after_set[31];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[32] <= 0;
    end
    else begin
      regs[32] <= after_set[32];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[33] <= 0;
    end
    else begin
      regs[33] <= after_set[33];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[34] <= 0;
    end
    else begin
      regs[34] <= after_set[34];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[35] <= 0;
    end
    else begin
      regs[35] <= after_set[35];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[36] <= 0;
    end
    else begin
      regs[36] <= after_set[36];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[37] <= 0;
    end
    else begin
      regs[37] <= after_set[37];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[38] <= 0;
    end
    else begin
      regs[38] <= after_set[38];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[39] <= 0;
    end
    else begin
      regs[39] <= after_set[39];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[40] <= 0;
    end
    else begin
      regs[40] <= after_set[40];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[41] <= 0;
    end
    else begin
      regs[41] <= after_set[41];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[42] <= 0;
    end
    else begin
      regs[42] <= after_set[42];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[43] <= 0;
    end
    else begin
      regs[43] <= after_set[43];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[44] <= 0;
    end
    else begin
      regs[44] <= after_set[44];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[45] <= 0;
    end
    else begin
      regs[45] <= after_set[45];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[46] <= 0;
    end
    else begin
      regs[46] <= after_set[46];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[47] <= 0;
    end
    else begin
      regs[47] <= after_set[47];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[48] <= 0;
    end
    else begin
      regs[48] <= after_set[48];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[49] <= 0;
    end
    else begin
      regs[49] <= after_set[49];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[50] <= 0;
    end
    else begin
      regs[50] <= after_set[50];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[51] <= 0;
    end
    else begin
      regs[51] <= after_set[51];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[52] <= 0;
    end
    else begin
      regs[52] <= after_set[52];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[53] <= 0;
    end
    else begin
      regs[53] <= after_set[53];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[54] <= 0;
    end
    else begin
      regs[54] <= after_set[54];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[55] <= 0;
    end
    else begin
      regs[55] <= after_set[55];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[56] <= 0;
    end
    else begin
      regs[56] <= after_set[56];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[57] <= 0;
    end
    else begin
      regs[57] <= after_set[57];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[58] <= 0;
    end
    else begin
      regs[58] <= after_set[58];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[59] <= 0;
    end
    else begin
      regs[59] <= after_set[59];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[60] <= 0;
    end
    else begin
      regs[60] <= after_set[60];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[61] <= 0;
    end
    else begin
      regs[61] <= after_set[61];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(reg_i=reg_i, value=reset_values[reg_i]):
  //         if s.reset:
  //           s.regs[reg_i].n = value
  //         else:
  //           s.regs[reg_i].n = s.after_set[reg_i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      regs[62] <= 0;
    end
    else begin
      regs[62] <= after_set[62];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 0))) begin
      write_inc[0] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[0] = regs[0];
      end
      else begin
        write_inc[0] = write_inc[-63];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[0] = write_inc[0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[0] = set_in_[0];
    end
    else begin
      after_set[0] = after_write[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 1))) begin
      write_inc[1] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[1] = regs[1];
      end
      else begin
        write_inc[1] = write_inc[-62];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[1] = write_inc[1];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[1] = set_in_[1];
    end
    else begin
      after_set[1] = after_write[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 2))) begin
      write_inc[2] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[2] = regs[2];
      end
      else begin
        write_inc[2] = write_inc[-61];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[2] = write_inc[2];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[2] = set_in_[2];
    end
    else begin
      after_set[2] = after_write[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 3))) begin
      write_inc[3] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[3] = regs[3];
      end
      else begin
        write_inc[3] = write_inc[-60];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[3] = write_inc[3];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[3] = set_in_[3];
    end
    else begin
      after_set[3] = after_write[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 4))) begin
      write_inc[4] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[4] = regs[4];
      end
      else begin
        write_inc[4] = write_inc[-59];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[4] = write_inc[4];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[4] = set_in_[4];
    end
    else begin
      after_set[4] = after_write[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 5))) begin
      write_inc[5] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[5] = regs[5];
      end
      else begin
        write_inc[5] = write_inc[-58];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[5] = write_inc[5];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[5] = set_in_[5];
    end
    else begin
      after_set[5] = after_write[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 6))) begin
      write_inc[6] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[6] = regs[6];
      end
      else begin
        write_inc[6] = write_inc[-57];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[6] = write_inc[6];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[6] = set_in_[6];
    end
    else begin
      after_set[6] = after_write[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 7))) begin
      write_inc[7] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[7] = regs[7];
      end
      else begin
        write_inc[7] = write_inc[-56];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[7] = write_inc[7];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[7] = set_in_[7];
    end
    else begin
      after_set[7] = after_write[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 8))) begin
      write_inc[8] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[8] = regs[8];
      end
      else begin
        write_inc[8] = write_inc[-55];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[8] = write_inc[8];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[8] = set_in_[8];
    end
    else begin
      after_set[8] = after_write[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 9))) begin
      write_inc[9] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[9] = regs[9];
      end
      else begin
        write_inc[9] = write_inc[-54];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[9] = write_inc[9];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[9] = set_in_[9];
    end
    else begin
      after_set[9] = after_write[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 10))) begin
      write_inc[10] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[10] = regs[10];
      end
      else begin
        write_inc[10] = write_inc[-53];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[10] = write_inc[10];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[10] = set_in_[10];
    end
    else begin
      after_set[10] = after_write[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 11))) begin
      write_inc[11] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[11] = regs[11];
      end
      else begin
        write_inc[11] = write_inc[-52];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[11] = write_inc[11];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[11] = set_in_[11];
    end
    else begin
      after_set[11] = after_write[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 12))) begin
      write_inc[12] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[12] = regs[12];
      end
      else begin
        write_inc[12] = write_inc[-51];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[12] = write_inc[12];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[12] = set_in_[12];
    end
    else begin
      after_set[12] = after_write[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 13))) begin
      write_inc[13] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[13] = regs[13];
      end
      else begin
        write_inc[13] = write_inc[-50];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[13] = write_inc[13];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[13] = set_in_[13];
    end
    else begin
      after_set[13] = after_write[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 14))) begin
      write_inc[14] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[14] = regs[14];
      end
      else begin
        write_inc[14] = write_inc[-49];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[14] = write_inc[14];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[14] = set_in_[14];
    end
    else begin
      after_set[14] = after_write[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 15))) begin
      write_inc[15] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[15] = regs[15];
      end
      else begin
        write_inc[15] = write_inc[-48];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[15] = write_inc[15];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[15] = set_in_[15];
    end
    else begin
      after_set[15] = after_write[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 16))) begin
      write_inc[16] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[16] = regs[16];
      end
      else begin
        write_inc[16] = write_inc[-47];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[16] = write_inc[16];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[16] = set_in_[16];
    end
    else begin
      after_set[16] = after_write[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 17))) begin
      write_inc[17] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[17] = regs[17];
      end
      else begin
        write_inc[17] = write_inc[-46];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[17] = write_inc[17];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[17] = set_in_[17];
    end
    else begin
      after_set[17] = after_write[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 18))) begin
      write_inc[18] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[18] = regs[18];
      end
      else begin
        write_inc[18] = write_inc[-45];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[18] = write_inc[18];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[18] = set_in_[18];
    end
    else begin
      after_set[18] = after_write[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 19))) begin
      write_inc[19] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[19] = regs[19];
      end
      else begin
        write_inc[19] = write_inc[-44];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[19] = write_inc[19];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[19] = set_in_[19];
    end
    else begin
      after_set[19] = after_write[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 20))) begin
      write_inc[20] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[20] = regs[20];
      end
      else begin
        write_inc[20] = write_inc[-43];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[20] = write_inc[20];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[20] = set_in_[20];
    end
    else begin
      after_set[20] = after_write[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 21))) begin
      write_inc[21] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[21] = regs[21];
      end
      else begin
        write_inc[21] = write_inc[-42];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[21] = write_inc[21];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[21] = set_in_[21];
    end
    else begin
      after_set[21] = after_write[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 22))) begin
      write_inc[22] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[22] = regs[22];
      end
      else begin
        write_inc[22] = write_inc[-41];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[22] = write_inc[22];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[22] = set_in_[22];
    end
    else begin
      after_set[22] = after_write[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 23))) begin
      write_inc[23] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[23] = regs[23];
      end
      else begin
        write_inc[23] = write_inc[-40];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[23] = write_inc[23];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[23] = set_in_[23];
    end
    else begin
      after_set[23] = after_write[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 24))) begin
      write_inc[24] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[24] = regs[24];
      end
      else begin
        write_inc[24] = write_inc[-39];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[24] = write_inc[24];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[24] = set_in_[24];
    end
    else begin
      after_set[24] = after_write[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 25))) begin
      write_inc[25] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[25] = regs[25];
      end
      else begin
        write_inc[25] = write_inc[-38];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[25] = write_inc[25];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[25] = set_in_[25];
    end
    else begin
      after_set[25] = after_write[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 26))) begin
      write_inc[26] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[26] = regs[26];
      end
      else begin
        write_inc[26] = write_inc[-37];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[26] = write_inc[26];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[26] = set_in_[26];
    end
    else begin
      after_set[26] = after_write[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 27))) begin
      write_inc[27] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[27] = regs[27];
      end
      else begin
        write_inc[27] = write_inc[-36];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[27] = write_inc[27];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[27] = set_in_[27];
    end
    else begin
      after_set[27] = after_write[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 28))) begin
      write_inc[28] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[28] = regs[28];
      end
      else begin
        write_inc[28] = write_inc[-35];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[28] = write_inc[28];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[28] = set_in_[28];
    end
    else begin
      after_set[28] = after_write[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 29))) begin
      write_inc[29] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[29] = regs[29];
      end
      else begin
        write_inc[29] = write_inc[-34];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[29] = write_inc[29];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[29] = set_in_[29];
    end
    else begin
      after_set[29] = after_write[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 30))) begin
      write_inc[30] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[30] = regs[30];
      end
      else begin
        write_inc[30] = write_inc[-33];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[30] = write_inc[30];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[30] = set_in_[30];
    end
    else begin
      after_set[30] = after_write[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 31))) begin
      write_inc[31] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[31] = regs[31];
      end
      else begin
        write_inc[31] = write_inc[-32];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[31] = write_inc[31];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[31] = set_in_[31];
    end
    else begin
      after_set[31] = after_write[31];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 32))) begin
      write_inc[32] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[32] = regs[32];
      end
      else begin
        write_inc[32] = write_inc[-31];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[32] = write_inc[32];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[32] = set_in_[32];
    end
    else begin
      after_set[32] = after_write[32];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 33))) begin
      write_inc[33] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[33] = regs[33];
      end
      else begin
        write_inc[33] = write_inc[-30];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[33] = write_inc[33];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[33] = set_in_[33];
    end
    else begin
      after_set[33] = after_write[33];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 34))) begin
      write_inc[34] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[34] = regs[34];
      end
      else begin
        write_inc[34] = write_inc[-29];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[34] = write_inc[34];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[34] = set_in_[34];
    end
    else begin
      after_set[34] = after_write[34];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 35))) begin
      write_inc[35] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[35] = regs[35];
      end
      else begin
        write_inc[35] = write_inc[-28];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[35] = write_inc[35];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[35] = set_in_[35];
    end
    else begin
      after_set[35] = after_write[35];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 36))) begin
      write_inc[36] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[36] = regs[36];
      end
      else begin
        write_inc[36] = write_inc[-27];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[36] = write_inc[36];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[36] = set_in_[36];
    end
    else begin
      after_set[36] = after_write[36];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 37))) begin
      write_inc[37] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[37] = regs[37];
      end
      else begin
        write_inc[37] = write_inc[-26];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[37] = write_inc[37];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[37] = set_in_[37];
    end
    else begin
      after_set[37] = after_write[37];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 38))) begin
      write_inc[38] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[38] = regs[38];
      end
      else begin
        write_inc[38] = write_inc[-25];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[38] = write_inc[38];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[38] = set_in_[38];
    end
    else begin
      after_set[38] = after_write[38];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 39))) begin
      write_inc[39] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[39] = regs[39];
      end
      else begin
        write_inc[39] = write_inc[-24];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[39] = write_inc[39];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[39] = set_in_[39];
    end
    else begin
      after_set[39] = after_write[39];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 40))) begin
      write_inc[40] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[40] = regs[40];
      end
      else begin
        write_inc[40] = write_inc[-23];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[40] = write_inc[40];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[40] = set_in_[40];
    end
    else begin
      after_set[40] = after_write[40];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 41))) begin
      write_inc[41] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[41] = regs[41];
      end
      else begin
        write_inc[41] = write_inc[-22];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[41] = write_inc[41];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[41] = set_in_[41];
    end
    else begin
      after_set[41] = after_write[41];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 42))) begin
      write_inc[42] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[42] = regs[42];
      end
      else begin
        write_inc[42] = write_inc[-21];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[42] = write_inc[42];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[42] = set_in_[42];
    end
    else begin
      after_set[42] = after_write[42];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 43))) begin
      write_inc[43] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[43] = regs[43];
      end
      else begin
        write_inc[43] = write_inc[-20];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[43] = write_inc[43];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[43] = set_in_[43];
    end
    else begin
      after_set[43] = after_write[43];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 44))) begin
      write_inc[44] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[44] = regs[44];
      end
      else begin
        write_inc[44] = write_inc[-19];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[44] = write_inc[44];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[44] = set_in_[44];
    end
    else begin
      after_set[44] = after_write[44];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 45))) begin
      write_inc[45] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[45] = regs[45];
      end
      else begin
        write_inc[45] = write_inc[-18];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[45] = write_inc[45];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[45] = set_in_[45];
    end
    else begin
      after_set[45] = after_write[45];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 46))) begin
      write_inc[46] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[46] = regs[46];
      end
      else begin
        write_inc[46] = write_inc[-17];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[46] = write_inc[46];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[46] = set_in_[46];
    end
    else begin
      after_set[46] = after_write[46];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 47))) begin
      write_inc[47] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[47] = regs[47];
      end
      else begin
        write_inc[47] = write_inc[-16];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[47] = write_inc[47];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[47] = set_in_[47];
    end
    else begin
      after_set[47] = after_write[47];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 48))) begin
      write_inc[48] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[48] = regs[48];
      end
      else begin
        write_inc[48] = write_inc[-15];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[48] = write_inc[48];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[48] = set_in_[48];
    end
    else begin
      after_set[48] = after_write[48];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 49))) begin
      write_inc[49] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[49] = regs[49];
      end
      else begin
        write_inc[49] = write_inc[-14];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[49] = write_inc[49];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[49] = set_in_[49];
    end
    else begin
      after_set[49] = after_write[49];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 50))) begin
      write_inc[50] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[50] = regs[50];
      end
      else begin
        write_inc[50] = write_inc[-13];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[50] = write_inc[50];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[50] = set_in_[50];
    end
    else begin
      after_set[50] = after_write[50];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 51))) begin
      write_inc[51] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[51] = regs[51];
      end
      else begin
        write_inc[51] = write_inc[-12];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[51] = write_inc[51];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[51] = set_in_[51];
    end
    else begin
      after_set[51] = after_write[51];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 52))) begin
      write_inc[52] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[52] = regs[52];
      end
      else begin
        write_inc[52] = write_inc[-11];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[52] = write_inc[52];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[52] = set_in_[52];
    end
    else begin
      after_set[52] = after_write[52];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 53))) begin
      write_inc[53] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[53] = regs[53];
      end
      else begin
        write_inc[53] = write_inc[-10];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[53] = write_inc[53];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[53] = set_in_[53];
    end
    else begin
      after_set[53] = after_write[53];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 54))) begin
      write_inc[54] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[54] = regs[54];
      end
      else begin
        write_inc[54] = write_inc[-9];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[54] = write_inc[54];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[54] = set_in_[54];
    end
    else begin
      after_set[54] = after_write[54];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 55))) begin
      write_inc[55] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[55] = regs[55];
      end
      else begin
        write_inc[55] = write_inc[-8];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[55] = write_inc[55];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[55] = set_in_[55];
    end
    else begin
      after_set[55] = after_write[55];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 56))) begin
      write_inc[56] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[56] = regs[56];
      end
      else begin
        write_inc[56] = write_inc[-7];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[56] = write_inc[56];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[56] = set_in_[56];
    end
    else begin
      after_set[56] = after_write[56];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 57))) begin
      write_inc[57] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[57] = regs[57];
      end
      else begin
        write_inc[57] = write_inc[-6];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[57] = write_inc[57];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[57] = set_in_[57];
    end
    else begin
      after_set[57] = after_write[57];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 58))) begin
      write_inc[58] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[58] = regs[58];
      end
      else begin
        write_inc[58] = write_inc[-5];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[58] = write_inc[58];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[58] = set_in_[58];
    end
    else begin
      after_set[58] = after_write[58];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 59))) begin
      write_inc[59] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[59] = regs[59];
      end
      else begin
        write_inc[59] = write_inc[-4];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[59] = write_inc[59];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[59] = set_in_[59];
    end
    else begin
      after_set[59] = after_write[59];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 60))) begin
      write_inc[60] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[60] = regs[60];
      end
      else begin
        write_inc[60] = write_inc[-3];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[60] = write_inc[60];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[60] = set_in_[60];
    end
    else begin
      after_set[60] = after_write[60];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 61))) begin
      write_inc[61] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[61] = regs[61];
      end
      else begin
        write_inc[61] = write_inc[-2];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[61] = write_inc[61];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[61] = set_in_[61];
    end
    else begin
      after_set[61] = after_write[61];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_write(reg_i=reg_i,
  //                          port=port,
  //                          i=port * nregs + reg_i,
  //                          j=(port - 1) * nregs + reg_i):
  //           if s.write_call[port] and s.write_addr[port] == reg_i:
  //             s.write_inc[i].v = s.write_data[port]
  //           elif port == 0:
  //             s.write_inc[i].v = s.regs[reg_i]
  //           else:
  //             s.write_inc[i].v = s.write_inc[j]

  // logic for handle_write()
  always @ (*) begin
    if ((write_call[0]&&(write_addr[0] == 62))) begin
      write_inc[62] = write_data[0];
    end
    else begin
      if ((0 == 0)) begin
        write_inc[62] = regs[62];
      end
      else begin
        write_inc[62] = write_inc[-1];
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_last(reg_i=reg_i, i=(num_write_ports - 1) * nregs + reg_i):
  //           s.after_write[reg_i].v = s.write_inc[i]

  // logic for update_last()
  always @ (*) begin
    after_write[62] = write_inc[62];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_set(reg_i=reg_i):
  //         if s.set_call:
  //           s.after_set[reg_i].v = s.set_in_[reg_i]
  //         else:
  //           s.after_set[reg_i].v = s.after_write[reg_i]

  // logic for handle_set()
  always @ (*) begin
    if (set_call) begin
      after_set[62] = set_in_[62];
    end
    else begin
      after_set[62] = after_write[62];
    end
  end


endmodule // RegisterFile_0x764ec1b6bf9dc34b

//-----------------------------------------------------------------------------
// Mux_0x7af68b5383bacfb2
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.mux {"dtype": 63, "nports": 2}
// PyMTL: verilator_xinit = zeros
module Mux_0x7af68b5383bacfb2
(
  input  logic [   0:0] clk,
  input  logic [  62:0] mux_in_$000,
  input  logic [  62:0] mux_in_$001,
  output logic  [  62:0] mux_out,
  input  logic [   0:0] mux_select,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nports = 2;


  // array declarations
  logic   [  62:0] mux_in_[0:1];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def select():
  //       assert s.mux_select < nports
  //       s.mux_out.v = s.mux_in_[s.mux_select]

  // logic for select()
  always @ (*) begin
    mux_out = mux_in_[mux_select];
  end


endmodule // Mux_0x7af68b5383bacfb2

//-----------------------------------------------------------------------------
// FreeList_0x2dd76b08b1ccb6ed
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.freelist {"free_alloc_bypass": false, "nslots": 63, "num_alloc_ports": 1, "num_free_ports": 2, "release_alloc_bypass": false, "used_slots_initial": 31}
// PyMTL: verilator_xinit = zeros
module FreeList_0x2dd76b08b1ccb6ed
(
  input  logic [   0:0] alloc_call$000,
  output logic [   5:0] alloc_index$000,
  output logic [  62:0] alloc_mask$000,
  output logic [   0:0] alloc_rdy$000,
  input  logic [   0:0] clk,
  input  logic [   0:0] free_call$000,
  input  logic [   0:0] free_call$001,
  input  logic [   5:0] free_index$000,
  input  logic [   5:0] free_index$001,
  input  logic [   0:0] release_call,
  input  logic [  62:0] release_mask,
  input  logic [   0:0] reset,
  input  logic [   0:0] set_call,
  input  logic [  62:0] set_state
);

  // logic declarations
  logic   [  62:0] free_masks$000;
  logic   [  62:0] free_masks$001;
  logic   [  62:0] free_masks$002;
  logic   [  62:0] alloc_inc$000;
  logic   [  62:0] alloc_inc$001;


  // register declarations
  logic    [  62:0] alloc_inc_base;
  logic    [  62:0] free_next;
  logic    [  62:0] free_next_base;
  logic    [  62:0] free_vector;

  // localparam declarations
  localparam num_alloc_ports = 1;
  localparam num_free_ports = 2;

  // free_encoders$000 temporaries
  logic   [   0:0] free_encoders$000$clk;
  logic   [   0:0] free_encoders$000$reset;
  logic   [   5:0] free_encoders$000$encode_number;
  logic   [  62:0] free_encoders$000$encode_onehot;

  OneHotEncoder_0x610bc488d4ab0a9b free_encoders$000
  (
    .clk           ( free_encoders$000$clk ),
    .reset         ( free_encoders$000$reset ),
    .encode_number ( free_encoders$000$encode_number ),
    .encode_onehot ( free_encoders$000$encode_onehot )
  );

  // free_encoders$001 temporaries
  logic   [   0:0] free_encoders$001$clk;
  logic   [   0:0] free_encoders$001$reset;
  logic   [   5:0] free_encoders$001$encode_number;
  logic   [  62:0] free_encoders$001$encode_onehot;

  OneHotEncoder_0x610bc488d4ab0a9b free_encoders$001
  (
    .clk           ( free_encoders$001$clk ),
    .reset         ( free_encoders$001$reset ),
    .encode_number ( free_encoders$001$encode_number ),
    .encode_onehot ( free_encoders$001$encode_onehot )
  );

  // alloc_decoders$000 temporaries
  logic   [   0:0] alloc_decoders$000$clk;
  logic   [   0:0] alloc_decoders$000$reset;
  logic   [  62:0] alloc_decoders$000$decode_signal;
  logic   [   0:0] alloc_decoders$000$decode_valid;
  logic   [   5:0] alloc_decoders$000$decode_decoded;

  PriorityDecoder_0x2e5c0266b41857fd alloc_decoders$000
  (
    .clk            ( alloc_decoders$000$clk ),
    .reset          ( alloc_decoders$000$reset ),
    .decode_signal  ( alloc_decoders$000$decode_signal ),
    .decode_valid   ( alloc_decoders$000$decode_valid ),
    .decode_decoded ( alloc_decoders$000$decode_decoded )
  );

  // alloc_encoders$000 temporaries
  logic   [   0:0] alloc_encoders$000$clk;
  logic   [   0:0] alloc_encoders$000$reset;
  logic   [   5:0] alloc_encoders$000$encode_number;
  logic   [  62:0] alloc_encoders$000$encode_onehot;

  OneHotEncoder_0x610bc488d4ab0a9b alloc_encoders$000
  (
    .clk           ( alloc_encoders$000$clk ),
    .reset         ( alloc_encoders$000$reset ),
    .encode_number ( alloc_encoders$000$encode_number ),
    .encode_onehot ( alloc_encoders$000$encode_onehot )
  );

  // set_mux temporaries
  logic   [  62:0] set_mux$mux_in_$000;
  logic   [  62:0] set_mux$mux_in_$001;
  logic   [   0:0] set_mux$clk;
  logic   [   0:0] set_mux$reset;
  logic   [   0:0] set_mux$mux_select;
  logic   [  62:0] set_mux$mux_out;

  Mux_0x7af68b5383bacfb2 set_mux
  (
    .mux_in_$000 ( set_mux$mux_in_$000 ),
    .mux_in_$001 ( set_mux$mux_in_$001 ),
    .clk         ( set_mux$clk ),
    .reset       ( set_mux$reset ),
    .mux_select  ( set_mux$mux_select ),
    .mux_out     ( set_mux$mux_out )
  );

  // signal connections
  assign alloc_decoders$000$clk           = clk;
  assign alloc_decoders$000$decode_signal = alloc_inc$000;
  assign alloc_decoders$000$reset         = reset;
  assign alloc_encoders$000$clk           = clk;
  assign alloc_encoders$000$encode_number = alloc_decoders$000$decode_decoded;
  assign alloc_encoders$000$reset         = reset;
  assign alloc_index$000                  = alloc_decoders$000$decode_decoded;
  assign alloc_mask$000                   = alloc_encoders$000$encode_onehot;
  assign alloc_rdy$000                    = alloc_decoders$000$decode_valid;
  assign free_encoders$000$clk            = clk;
  assign free_encoders$000$encode_number  = free_index$000;
  assign free_encoders$000$reset          = reset;
  assign free_encoders$001$clk            = clk;
  assign free_encoders$001$encode_number  = free_index$001;
  assign free_encoders$001$reset          = reset;
  assign free_masks$000                   = 63'd0;
  assign set_mux$clk                      = clk;
  assign set_mux$mux_in_$000              = free_next;
  assign set_mux$mux_in_$001              = set_state;
  assign set_mux$mux_select               = set_call;
  assign set_mux$reset                    = reset;

  // array declarations
  logic   [   0:0] alloc_call[0:0];
  assign alloc_call[  0] = alloc_call$000;
  logic   [  62:0] alloc_encoders$encode_onehot[0:0];
  assign alloc_encoders$encode_onehot[  0] = alloc_encoders$000$encode_onehot;
  logic    [  62:0] alloc_inc[0:1];
  assign alloc_inc$000 = alloc_inc[  0];
  assign alloc_inc$001 = alloc_inc[  1];
  logic   [   0:0] free_call[0:1];
  assign free_call[  0] = free_call$000;
  assign free_call[  1] = free_call$001;
  logic   [  62:0] free_encoders$encode_onehot[0:1];
  assign free_encoders$encode_onehot[  0] = free_encoders$000$encode_onehot;
  assign free_encoders$encode_onehot[  1] = free_encoders$001$encode_onehot;
  logic    [  62:0] free_masks[0:2];
  assign free_masks$000 = free_masks[  0];
  assign free_masks$001 = free_masks[  1];
  assign free_masks$002 = free_masks[  2];

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[0] <= 0;
    end
    else begin
      free_vector[0] <= set_mux$mux_out[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[1] <= 0;
    end
    else begin
      free_vector[1] <= set_mux$mux_out[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[2] <= 0;
    end
    else begin
      free_vector[2] <= set_mux$mux_out[2];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[3] <= 0;
    end
    else begin
      free_vector[3] <= set_mux$mux_out[3];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[4] <= 0;
    end
    else begin
      free_vector[4] <= set_mux$mux_out[4];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[5] <= 0;
    end
    else begin
      free_vector[5] <= set_mux$mux_out[5];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[6] <= 0;
    end
    else begin
      free_vector[6] <= set_mux$mux_out[6];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[7] <= 0;
    end
    else begin
      free_vector[7] <= set_mux$mux_out[7];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[8] <= 0;
    end
    else begin
      free_vector[8] <= set_mux$mux_out[8];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[9] <= 0;
    end
    else begin
      free_vector[9] <= set_mux$mux_out[9];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[10] <= 0;
    end
    else begin
      free_vector[10] <= set_mux$mux_out[10];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[11] <= 0;
    end
    else begin
      free_vector[11] <= set_mux$mux_out[11];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[12] <= 0;
    end
    else begin
      free_vector[12] <= set_mux$mux_out[12];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[13] <= 0;
    end
    else begin
      free_vector[13] <= set_mux$mux_out[13];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[14] <= 0;
    end
    else begin
      free_vector[14] <= set_mux$mux_out[14];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[15] <= 0;
    end
    else begin
      free_vector[15] <= set_mux$mux_out[15];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[16] <= 0;
    end
    else begin
      free_vector[16] <= set_mux$mux_out[16];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[17] <= 0;
    end
    else begin
      free_vector[17] <= set_mux$mux_out[17];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[18] <= 0;
    end
    else begin
      free_vector[18] <= set_mux$mux_out[18];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[19] <= 0;
    end
    else begin
      free_vector[19] <= set_mux$mux_out[19];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[20] <= 0;
    end
    else begin
      free_vector[20] <= set_mux$mux_out[20];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[21] <= 0;
    end
    else begin
      free_vector[21] <= set_mux$mux_out[21];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[22] <= 0;
    end
    else begin
      free_vector[22] <= set_mux$mux_out[22];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[23] <= 0;
    end
    else begin
      free_vector[23] <= set_mux$mux_out[23];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[24] <= 0;
    end
    else begin
      free_vector[24] <= set_mux$mux_out[24];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[25] <= 0;
    end
    else begin
      free_vector[25] <= set_mux$mux_out[25];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[26] <= 0;
    end
    else begin
      free_vector[26] <= set_mux$mux_out[26];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[27] <= 0;
    end
    else begin
      free_vector[27] <= set_mux$mux_out[27];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[28] <= 0;
    end
    else begin
      free_vector[28] <= set_mux$mux_out[28];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[29] <= 0;
    end
    else begin
      free_vector[29] <= set_mux$mux_out[29];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[30] <= 0;
    end
    else begin
      free_vector[30] <= set_mux$mux_out[30];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[31] <= 1;
    end
    else begin
      free_vector[31] <= set_mux$mux_out[31];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[32] <= 1;
    end
    else begin
      free_vector[32] <= set_mux$mux_out[32];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[33] <= 1;
    end
    else begin
      free_vector[33] <= set_mux$mux_out[33];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[34] <= 1;
    end
    else begin
      free_vector[34] <= set_mux$mux_out[34];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[35] <= 1;
    end
    else begin
      free_vector[35] <= set_mux$mux_out[35];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[36] <= 1;
    end
    else begin
      free_vector[36] <= set_mux$mux_out[36];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[37] <= 1;
    end
    else begin
      free_vector[37] <= set_mux$mux_out[37];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[38] <= 1;
    end
    else begin
      free_vector[38] <= set_mux$mux_out[38];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[39] <= 1;
    end
    else begin
      free_vector[39] <= set_mux$mux_out[39];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[40] <= 1;
    end
    else begin
      free_vector[40] <= set_mux$mux_out[40];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[41] <= 1;
    end
    else begin
      free_vector[41] <= set_mux$mux_out[41];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[42] <= 1;
    end
    else begin
      free_vector[42] <= set_mux$mux_out[42];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[43] <= 1;
    end
    else begin
      free_vector[43] <= set_mux$mux_out[43];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[44] <= 1;
    end
    else begin
      free_vector[44] <= set_mux$mux_out[44];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[45] <= 1;
    end
    else begin
      free_vector[45] <= set_mux$mux_out[45];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[46] <= 1;
    end
    else begin
      free_vector[46] <= set_mux$mux_out[46];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[47] <= 1;
    end
    else begin
      free_vector[47] <= set_mux$mux_out[47];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[48] <= 1;
    end
    else begin
      free_vector[48] <= set_mux$mux_out[48];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[49] <= 1;
    end
    else begin
      free_vector[49] <= set_mux$mux_out[49];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[50] <= 1;
    end
    else begin
      free_vector[50] <= set_mux$mux_out[50];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[51] <= 1;
    end
    else begin
      free_vector[51] <= set_mux$mux_out[51];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[52] <= 1;
    end
    else begin
      free_vector[52] <= set_mux$mux_out[52];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[53] <= 1;
    end
    else begin
      free_vector[53] <= set_mux$mux_out[53];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[54] <= 1;
    end
    else begin
      free_vector[54] <= set_mux$mux_out[54];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[55] <= 1;
    end
    else begin
      free_vector[55] <= set_mux$mux_out[55];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[56] <= 1;
    end
    else begin
      free_vector[56] <= set_mux$mux_out[56];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[57] <= 1;
    end
    else begin
      free_vector[57] <= set_mux$mux_out[57];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[58] <= 1;
    end
    else begin
      free_vector[58] <= set_mux$mux_out[58];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[59] <= 1;
    end
    else begin
      free_vector[59] <= set_mux$mux_out[59];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[60] <= 1;
    end
    else begin
      free_vector[60] <= set_mux$mux_out[60];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[61] <= 1;
    end
    else begin
      free_vector[61] <= set_mux$mux_out[61];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update(i=i, free=(1 if i >= used_slots_initial else 0)):
  //         if s.reset:
  //           s.free_vector[i].n = free
  //         else:
  //           s.free_vector[i].n = s.set_mux.mux_out[i]

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      free_vector[62] <= 1;
    end
    else begin
      free_vector[62] <= set_mux$mux_out[62];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_free(n=i + 1, i=i):
  //         if s.free_call[i]:
  //           s.free_masks[n].v = s.free_masks[i] | s.free_encoders[i].encode_onehot
  //         else:
  //           s.free_masks[n].v = s.free_masks[i]

  // logic for handle_free()
  always @ (*) begin
    if (free_call[0]) begin
      free_masks[1] = (free_masks[0]|free_encoders$encode_onehot[0]);
    end
    else begin
      free_masks[1] = free_masks[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_free(n=i + 1, i=i):
  //         if s.free_call[i]:
  //           s.free_masks[n].v = s.free_masks[i] | s.free_encoders[i].encode_onehot
  //         else:
  //           s.free_masks[n].v = s.free_masks[i]

  // logic for handle_free()
  always @ (*) begin
    if (free_call[1]) begin
      free_masks[2] = (free_masks[1]|free_encoders$encode_onehot[1]);
    end
    else begin
      free_masks[2] = free_masks[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_alloc_inc_base():
  //         s.alloc_inc_base.v = s.free_vector

  // logic for compute_alloc_inc_base()
  always @ (*) begin
    alloc_inc_base = free_vector;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_alloc_inc_0():
  //         s.alloc_inc[0].v = s.alloc_inc_base

  // logic for compute_alloc_inc_0()
  always @ (*) begin
    alloc_inc[0] = alloc_inc_base;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_alloc(n=i + 1, i=i):
  //         if s.alloc_call[i]:
  //           s.alloc_inc[n].v = s.alloc_inc[i] & (
  //               ~s.alloc_encoders[i].encode_onehot)
  //         else:
  //           s.alloc_inc[n].v = s.alloc_inc[i]

  // logic for handle_alloc()
  always @ (*) begin
    if (alloc_call[0]) begin
      alloc_inc[1] = (alloc_inc[0]&~alloc_encoders$encode_onehot[0]);
    end
    else begin
      alloc_inc[1] = alloc_inc[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_free_next_base():
  //         if s.release_call:
  //           s.free_next_base.v = s.alloc_inc[num_alloc_ports] | s.release_mask
  //         else:
  //           s.free_next_base.v = s.alloc_inc[num_alloc_ports]

  // logic for compute_free_next_base()
  always @ (*) begin
    if (release_call) begin
      free_next_base = (alloc_inc[num_alloc_ports]|release_mask);
    end
    else begin
      free_next_base = alloc_inc[num_alloc_ports];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_free():
  //         s.free_next.v = s.free_next_base | s.free_masks[num_free_ports]

  // logic for compute_free()
  always @ (*) begin
    free_next = (free_next_base|free_masks[num_free_ports]);
  end


endmodule // FreeList_0x2dd76b08b1ccb6ed

//-----------------------------------------------------------------------------
// OneHotEncoder_0x610bc488d4ab0a9b
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.onehot {"enable": false, "noutbits": 63}
// PyMTL: verilator_xinit = zeros
module OneHotEncoder_0x610bc488d4ab0a9b
(
  input  logic [   0:0] clk,
  input  logic [   5:0] encode_number,
  output logic  [  62:0] encode_onehot,
  input  logic [   0:0] reset
);



  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[0] = (encode_number == 0);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[1] = (encode_number == 1);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[2] = (encode_number == 2);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[3] = (encode_number == 3);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[4] = (encode_number == 4);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[5] = (encode_number == 5);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[6] = (encode_number == 6);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[7] = (encode_number == 7);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[8] = (encode_number == 8);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[9] = (encode_number == 9);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[10] = (encode_number == 10);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[11] = (encode_number == 11);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[12] = (encode_number == 12);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[13] = (encode_number == 13);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[14] = (encode_number == 14);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[15] = (encode_number == 15);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[16] = (encode_number == 16);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[17] = (encode_number == 17);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[18] = (encode_number == 18);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[19] = (encode_number == 19);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[20] = (encode_number == 20);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[21] = (encode_number == 21);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[22] = (encode_number == 22);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[23] = (encode_number == 23);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[24] = (encode_number == 24);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[25] = (encode_number == 25);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[26] = (encode_number == 26);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[27] = (encode_number == 27);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[28] = (encode_number == 28);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[29] = (encode_number == 29);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[30] = (encode_number == 30);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[31] = (encode_number == 31);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[32] = (encode_number == 32);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[33] = (encode_number == 33);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[34] = (encode_number == 34);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[35] = (encode_number == 35);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[36] = (encode_number == 36);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[37] = (encode_number == 37);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[38] = (encode_number == 38);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[39] = (encode_number == 39);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[40] = (encode_number == 40);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[41] = (encode_number == 41);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[42] = (encode_number == 42);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[43] = (encode_number == 43);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[44] = (encode_number == 44);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[45] = (encode_number == 45);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[46] = (encode_number == 46);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[47] = (encode_number == 47);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[48] = (encode_number == 48);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[49] = (encode_number == 49);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[50] = (encode_number == 50);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[51] = (encode_number == 51);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[52] = (encode_number == 52);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[53] = (encode_number == 53);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[54] = (encode_number == 54);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[55] = (encode_number == 55);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[56] = (encode_number == 56);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[57] = (encode_number == 57);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[58] = (encode_number == 58);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[59] = (encode_number == 59);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[60] = (encode_number == 60);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[61] = (encode_number == 61);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[62] = (encode_number == 62);
  end


endmodule // OneHotEncoder_0x610bc488d4ab0a9b

//-----------------------------------------------------------------------------
// PriorityDecoder_0x2e5c0266b41857fd
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.coders {"inwidth": 63}
// PyMTL: verilator_xinit = zeros
module PriorityDecoder_0x2e5c0266b41857fd
(
  input  logic [   0:0] clk,
  output logic [   5:0] decode_decoded,
  input  logic [  62:0] decode_signal,
  output logic [   0:0] decode_valid,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   5:0] outs$000;
  logic   [   5:0] outs$001;
  logic   [   5:0] outs$002;
  logic   [   5:0] outs$003;
  logic   [   5:0] outs$004;
  logic   [   5:0] outs$005;
  logic   [   5:0] outs$006;
  logic   [   5:0] outs$007;
  logic   [   5:0] outs$008;
  logic   [   5:0] outs$009;
  logic   [   5:0] outs$010;
  logic   [   5:0] outs$011;
  logic   [   5:0] outs$012;
  logic   [   5:0] outs$013;
  logic   [   5:0] outs$014;
  logic   [   5:0] outs$015;
  logic   [   5:0] outs$016;
  logic   [   5:0] outs$017;
  logic   [   5:0] outs$018;
  logic   [   5:0] outs$019;
  logic   [   5:0] outs$020;
  logic   [   5:0] outs$021;
  logic   [   5:0] outs$022;
  logic   [   5:0] outs$023;
  logic   [   5:0] outs$024;
  logic   [   5:0] outs$025;
  logic   [   5:0] outs$026;
  logic   [   5:0] outs$027;
  logic   [   5:0] outs$028;
  logic   [   5:0] outs$029;
  logic   [   5:0] outs$030;
  logic   [   5:0] outs$031;
  logic   [   5:0] outs$032;
  logic   [   5:0] outs$033;
  logic   [   5:0] outs$034;
  logic   [   5:0] outs$035;
  logic   [   5:0] outs$036;
  logic   [   5:0] outs$037;
  logic   [   5:0] outs$038;
  logic   [   5:0] outs$039;
  logic   [   5:0] outs$040;
  logic   [   5:0] outs$041;
  logic   [   5:0] outs$042;
  logic   [   5:0] outs$043;
  logic   [   5:0] outs$044;
  logic   [   5:0] outs$045;
  logic   [   5:0] outs$046;
  logic   [   5:0] outs$047;
  logic   [   5:0] outs$048;
  logic   [   5:0] outs$049;
  logic   [   5:0] outs$050;
  logic   [   5:0] outs$051;
  logic   [   5:0] outs$052;
  logic   [   5:0] outs$053;
  logic   [   5:0] outs$054;
  logic   [   5:0] outs$055;
  logic   [   5:0] outs$056;
  logic   [   5:0] outs$057;
  logic   [   5:0] outs$058;
  logic   [   5:0] outs$059;
  logic   [   5:0] outs$060;
  logic   [   5:0] outs$061;
  logic   [   5:0] outs$062;
  logic   [   5:0] outs$063;
  logic   [   0:0] valid$000;
  logic   [   0:0] valid$001;
  logic   [   0:0] valid$002;
  logic   [   0:0] valid$003;
  logic   [   0:0] valid$004;
  logic   [   0:0] valid$005;
  logic   [   0:0] valid$006;
  logic   [   0:0] valid$007;
  logic   [   0:0] valid$008;
  logic   [   0:0] valid$009;
  logic   [   0:0] valid$010;
  logic   [   0:0] valid$011;
  logic   [   0:0] valid$012;
  logic   [   0:0] valid$013;
  logic   [   0:0] valid$014;
  logic   [   0:0] valid$015;
  logic   [   0:0] valid$016;
  logic   [   0:0] valid$017;
  logic   [   0:0] valid$018;
  logic   [   0:0] valid$019;
  logic   [   0:0] valid$020;
  logic   [   0:0] valid$021;
  logic   [   0:0] valid$022;
  logic   [   0:0] valid$023;
  logic   [   0:0] valid$024;
  logic   [   0:0] valid$025;
  logic   [   0:0] valid$026;
  logic   [   0:0] valid$027;
  logic   [   0:0] valid$028;
  logic   [   0:0] valid$029;
  logic   [   0:0] valid$030;
  logic   [   0:0] valid$031;
  logic   [   0:0] valid$032;
  logic   [   0:0] valid$033;
  logic   [   0:0] valid$034;
  logic   [   0:0] valid$035;
  logic   [   0:0] valid$036;
  logic   [   0:0] valid$037;
  logic   [   0:0] valid$038;
  logic   [   0:0] valid$039;
  logic   [   0:0] valid$040;
  logic   [   0:0] valid$041;
  logic   [   0:0] valid$042;
  logic   [   0:0] valid$043;
  logic   [   0:0] valid$044;
  logic   [   0:0] valid$045;
  logic   [   0:0] valid$046;
  logic   [   0:0] valid$047;
  logic   [   0:0] valid$048;
  logic   [   0:0] valid$049;
  logic   [   0:0] valid$050;
  logic   [   0:0] valid$051;
  logic   [   0:0] valid$052;
  logic   [   0:0] valid$053;
  logic   [   0:0] valid$054;
  logic   [   0:0] valid$055;
  logic   [   0:0] valid$056;
  logic   [   0:0] valid$057;
  logic   [   0:0] valid$058;
  logic   [   0:0] valid$059;
  logic   [   0:0] valid$060;
  logic   [   0:0] valid$061;
  logic   [   0:0] valid$062;
  logic   [   0:0] valid$063;


  // signal connections
  assign decode_decoded = outs$063;
  assign decode_valid   = valid$063;
  assign outs$000       = 6'd0;
  assign valid$000      = 1'd0;

  // array declarations
  logic    [   5:0] outs[0:63];
  assign outs$000 = outs[  0];
  assign outs$001 = outs[  1];
  assign outs$002 = outs[  2];
  assign outs$003 = outs[  3];
  assign outs$004 = outs[  4];
  assign outs$005 = outs[  5];
  assign outs$006 = outs[  6];
  assign outs$007 = outs[  7];
  assign outs$008 = outs[  8];
  assign outs$009 = outs[  9];
  assign outs$010 = outs[ 10];
  assign outs$011 = outs[ 11];
  assign outs$012 = outs[ 12];
  assign outs$013 = outs[ 13];
  assign outs$014 = outs[ 14];
  assign outs$015 = outs[ 15];
  assign outs$016 = outs[ 16];
  assign outs$017 = outs[ 17];
  assign outs$018 = outs[ 18];
  assign outs$019 = outs[ 19];
  assign outs$020 = outs[ 20];
  assign outs$021 = outs[ 21];
  assign outs$022 = outs[ 22];
  assign outs$023 = outs[ 23];
  assign outs$024 = outs[ 24];
  assign outs$025 = outs[ 25];
  assign outs$026 = outs[ 26];
  assign outs$027 = outs[ 27];
  assign outs$028 = outs[ 28];
  assign outs$029 = outs[ 29];
  assign outs$030 = outs[ 30];
  assign outs$031 = outs[ 31];
  assign outs$032 = outs[ 32];
  assign outs$033 = outs[ 33];
  assign outs$034 = outs[ 34];
  assign outs$035 = outs[ 35];
  assign outs$036 = outs[ 36];
  assign outs$037 = outs[ 37];
  assign outs$038 = outs[ 38];
  assign outs$039 = outs[ 39];
  assign outs$040 = outs[ 40];
  assign outs$041 = outs[ 41];
  assign outs$042 = outs[ 42];
  assign outs$043 = outs[ 43];
  assign outs$044 = outs[ 44];
  assign outs$045 = outs[ 45];
  assign outs$046 = outs[ 46];
  assign outs$047 = outs[ 47];
  assign outs$048 = outs[ 48];
  assign outs$049 = outs[ 49];
  assign outs$050 = outs[ 50];
  assign outs$051 = outs[ 51];
  assign outs$052 = outs[ 52];
  assign outs$053 = outs[ 53];
  assign outs$054 = outs[ 54];
  assign outs$055 = outs[ 55];
  assign outs$056 = outs[ 56];
  assign outs$057 = outs[ 57];
  assign outs$058 = outs[ 58];
  assign outs$059 = outs[ 59];
  assign outs$060 = outs[ 60];
  assign outs$061 = outs[ 61];
  assign outs$062 = outs[ 62];
  assign outs$063 = outs[ 63];
  logic    [   0:0] valid[0:63];
  assign valid$000 = valid[  0];
  assign valid$001 = valid[  1];
  assign valid$002 = valid[  2];
  assign valid$003 = valid[  3];
  assign valid$004 = valid[  4];
  assign valid$005 = valid[  5];
  assign valid$006 = valid[  6];
  assign valid$007 = valid[  7];
  assign valid$008 = valid[  8];
  assign valid$009 = valid[  9];
  assign valid$010 = valid[ 10];
  assign valid$011 = valid[ 11];
  assign valid$012 = valid[ 12];
  assign valid$013 = valid[ 13];
  assign valid$014 = valid[ 14];
  assign valid$015 = valid[ 15];
  assign valid$016 = valid[ 16];
  assign valid$017 = valid[ 17];
  assign valid$018 = valid[ 18];
  assign valid$019 = valid[ 19];
  assign valid$020 = valid[ 20];
  assign valid$021 = valid[ 21];
  assign valid$022 = valid[ 22];
  assign valid$023 = valid[ 23];
  assign valid$024 = valid[ 24];
  assign valid$025 = valid[ 25];
  assign valid$026 = valid[ 26];
  assign valid$027 = valid[ 27];
  assign valid$028 = valid[ 28];
  assign valid$029 = valid[ 29];
  assign valid$030 = valid[ 30];
  assign valid$031 = valid[ 31];
  assign valid$032 = valid[ 32];
  assign valid$033 = valid[ 33];
  assign valid$034 = valid[ 34];
  assign valid$035 = valid[ 35];
  assign valid$036 = valid[ 36];
  assign valid$037 = valid[ 37];
  assign valid$038 = valid[ 38];
  assign valid$039 = valid[ 39];
  assign valid$040 = valid[ 40];
  assign valid$041 = valid[ 41];
  assign valid$042 = valid[ 42];
  assign valid$043 = valid[ 43];
  assign valid$044 = valid[ 44];
  assign valid$045 = valid[ 45];
  assign valid$046 = valid[ 46];
  assign valid$047 = valid[ 47];
  assign valid$048 = valid[ 48];
  assign valid$049 = valid[ 49];
  assign valid$050 = valid[ 50];
  assign valid$051 = valid[ 51];
  assign valid$052 = valid[ 52];
  assign valid$053 = valid[ 53];
  assign valid$054 = valid[ 54];
  assign valid$055 = valid[ 55];
  assign valid$056 = valid[ 56];
  assign valid$057 = valid[ 57];
  assign valid$058 = valid[ 58];
  assign valid$059 = valid[ 59];
  assign valid$060 = valid[ 60];
  assign valid$061 = valid[ 61];
  assign valid$062 = valid[ 62];
  assign valid$063 = valid[ 63];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[0]) begin
      valid[1] = 1;
      outs[1] = outs[0];
    end
    else begin
      if (decode_signal[0]) begin
        valid[1] = 1;
        outs[1] = 0;
      end
      else begin
        valid[1] = 0;
        outs[1] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[1]) begin
      valid[2] = 1;
      outs[2] = outs[1];
    end
    else begin
      if (decode_signal[1]) begin
        valid[2] = 1;
        outs[2] = 1;
      end
      else begin
        valid[2] = 0;
        outs[2] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[2]) begin
      valid[3] = 1;
      outs[3] = outs[2];
    end
    else begin
      if (decode_signal[2]) begin
        valid[3] = 1;
        outs[3] = 2;
      end
      else begin
        valid[3] = 0;
        outs[3] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[3]) begin
      valid[4] = 1;
      outs[4] = outs[3];
    end
    else begin
      if (decode_signal[3]) begin
        valid[4] = 1;
        outs[4] = 3;
      end
      else begin
        valid[4] = 0;
        outs[4] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[4]) begin
      valid[5] = 1;
      outs[5] = outs[4];
    end
    else begin
      if (decode_signal[4]) begin
        valid[5] = 1;
        outs[5] = 4;
      end
      else begin
        valid[5] = 0;
        outs[5] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[5]) begin
      valid[6] = 1;
      outs[6] = outs[5];
    end
    else begin
      if (decode_signal[5]) begin
        valid[6] = 1;
        outs[6] = 5;
      end
      else begin
        valid[6] = 0;
        outs[6] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[6]) begin
      valid[7] = 1;
      outs[7] = outs[6];
    end
    else begin
      if (decode_signal[6]) begin
        valid[7] = 1;
        outs[7] = 6;
      end
      else begin
        valid[7] = 0;
        outs[7] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[7]) begin
      valid[8] = 1;
      outs[8] = outs[7];
    end
    else begin
      if (decode_signal[7]) begin
        valid[8] = 1;
        outs[8] = 7;
      end
      else begin
        valid[8] = 0;
        outs[8] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[8]) begin
      valid[9] = 1;
      outs[9] = outs[8];
    end
    else begin
      if (decode_signal[8]) begin
        valid[9] = 1;
        outs[9] = 8;
      end
      else begin
        valid[9] = 0;
        outs[9] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[9]) begin
      valid[10] = 1;
      outs[10] = outs[9];
    end
    else begin
      if (decode_signal[9]) begin
        valid[10] = 1;
        outs[10] = 9;
      end
      else begin
        valid[10] = 0;
        outs[10] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[10]) begin
      valid[11] = 1;
      outs[11] = outs[10];
    end
    else begin
      if (decode_signal[10]) begin
        valid[11] = 1;
        outs[11] = 10;
      end
      else begin
        valid[11] = 0;
        outs[11] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[11]) begin
      valid[12] = 1;
      outs[12] = outs[11];
    end
    else begin
      if (decode_signal[11]) begin
        valid[12] = 1;
        outs[12] = 11;
      end
      else begin
        valid[12] = 0;
        outs[12] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[12]) begin
      valid[13] = 1;
      outs[13] = outs[12];
    end
    else begin
      if (decode_signal[12]) begin
        valid[13] = 1;
        outs[13] = 12;
      end
      else begin
        valid[13] = 0;
        outs[13] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[13]) begin
      valid[14] = 1;
      outs[14] = outs[13];
    end
    else begin
      if (decode_signal[13]) begin
        valid[14] = 1;
        outs[14] = 13;
      end
      else begin
        valid[14] = 0;
        outs[14] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[14]) begin
      valid[15] = 1;
      outs[15] = outs[14];
    end
    else begin
      if (decode_signal[14]) begin
        valid[15] = 1;
        outs[15] = 14;
      end
      else begin
        valid[15] = 0;
        outs[15] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[15]) begin
      valid[16] = 1;
      outs[16] = outs[15];
    end
    else begin
      if (decode_signal[15]) begin
        valid[16] = 1;
        outs[16] = 15;
      end
      else begin
        valid[16] = 0;
        outs[16] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[16]) begin
      valid[17] = 1;
      outs[17] = outs[16];
    end
    else begin
      if (decode_signal[16]) begin
        valid[17] = 1;
        outs[17] = 16;
      end
      else begin
        valid[17] = 0;
        outs[17] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[17]) begin
      valid[18] = 1;
      outs[18] = outs[17];
    end
    else begin
      if (decode_signal[17]) begin
        valid[18] = 1;
        outs[18] = 17;
      end
      else begin
        valid[18] = 0;
        outs[18] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[18]) begin
      valid[19] = 1;
      outs[19] = outs[18];
    end
    else begin
      if (decode_signal[18]) begin
        valid[19] = 1;
        outs[19] = 18;
      end
      else begin
        valid[19] = 0;
        outs[19] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[19]) begin
      valid[20] = 1;
      outs[20] = outs[19];
    end
    else begin
      if (decode_signal[19]) begin
        valid[20] = 1;
        outs[20] = 19;
      end
      else begin
        valid[20] = 0;
        outs[20] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[20]) begin
      valid[21] = 1;
      outs[21] = outs[20];
    end
    else begin
      if (decode_signal[20]) begin
        valid[21] = 1;
        outs[21] = 20;
      end
      else begin
        valid[21] = 0;
        outs[21] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[21]) begin
      valid[22] = 1;
      outs[22] = outs[21];
    end
    else begin
      if (decode_signal[21]) begin
        valid[22] = 1;
        outs[22] = 21;
      end
      else begin
        valid[22] = 0;
        outs[22] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[22]) begin
      valid[23] = 1;
      outs[23] = outs[22];
    end
    else begin
      if (decode_signal[22]) begin
        valid[23] = 1;
        outs[23] = 22;
      end
      else begin
        valid[23] = 0;
        outs[23] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[23]) begin
      valid[24] = 1;
      outs[24] = outs[23];
    end
    else begin
      if (decode_signal[23]) begin
        valid[24] = 1;
        outs[24] = 23;
      end
      else begin
        valid[24] = 0;
        outs[24] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[24]) begin
      valid[25] = 1;
      outs[25] = outs[24];
    end
    else begin
      if (decode_signal[24]) begin
        valid[25] = 1;
        outs[25] = 24;
      end
      else begin
        valid[25] = 0;
        outs[25] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[25]) begin
      valid[26] = 1;
      outs[26] = outs[25];
    end
    else begin
      if (decode_signal[25]) begin
        valid[26] = 1;
        outs[26] = 25;
      end
      else begin
        valid[26] = 0;
        outs[26] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[26]) begin
      valid[27] = 1;
      outs[27] = outs[26];
    end
    else begin
      if (decode_signal[26]) begin
        valid[27] = 1;
        outs[27] = 26;
      end
      else begin
        valid[27] = 0;
        outs[27] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[27]) begin
      valid[28] = 1;
      outs[28] = outs[27];
    end
    else begin
      if (decode_signal[27]) begin
        valid[28] = 1;
        outs[28] = 27;
      end
      else begin
        valid[28] = 0;
        outs[28] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[28]) begin
      valid[29] = 1;
      outs[29] = outs[28];
    end
    else begin
      if (decode_signal[28]) begin
        valid[29] = 1;
        outs[29] = 28;
      end
      else begin
        valid[29] = 0;
        outs[29] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[29]) begin
      valid[30] = 1;
      outs[30] = outs[29];
    end
    else begin
      if (decode_signal[29]) begin
        valid[30] = 1;
        outs[30] = 29;
      end
      else begin
        valid[30] = 0;
        outs[30] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[30]) begin
      valid[31] = 1;
      outs[31] = outs[30];
    end
    else begin
      if (decode_signal[30]) begin
        valid[31] = 1;
        outs[31] = 30;
      end
      else begin
        valid[31] = 0;
        outs[31] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[31]) begin
      valid[32] = 1;
      outs[32] = outs[31];
    end
    else begin
      if (decode_signal[31]) begin
        valid[32] = 1;
        outs[32] = 31;
      end
      else begin
        valid[32] = 0;
        outs[32] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[32]) begin
      valid[33] = 1;
      outs[33] = outs[32];
    end
    else begin
      if (decode_signal[32]) begin
        valid[33] = 1;
        outs[33] = 32;
      end
      else begin
        valid[33] = 0;
        outs[33] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[33]) begin
      valid[34] = 1;
      outs[34] = outs[33];
    end
    else begin
      if (decode_signal[33]) begin
        valid[34] = 1;
        outs[34] = 33;
      end
      else begin
        valid[34] = 0;
        outs[34] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[34]) begin
      valid[35] = 1;
      outs[35] = outs[34];
    end
    else begin
      if (decode_signal[34]) begin
        valid[35] = 1;
        outs[35] = 34;
      end
      else begin
        valid[35] = 0;
        outs[35] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[35]) begin
      valid[36] = 1;
      outs[36] = outs[35];
    end
    else begin
      if (decode_signal[35]) begin
        valid[36] = 1;
        outs[36] = 35;
      end
      else begin
        valid[36] = 0;
        outs[36] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[36]) begin
      valid[37] = 1;
      outs[37] = outs[36];
    end
    else begin
      if (decode_signal[36]) begin
        valid[37] = 1;
        outs[37] = 36;
      end
      else begin
        valid[37] = 0;
        outs[37] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[37]) begin
      valid[38] = 1;
      outs[38] = outs[37];
    end
    else begin
      if (decode_signal[37]) begin
        valid[38] = 1;
        outs[38] = 37;
      end
      else begin
        valid[38] = 0;
        outs[38] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[38]) begin
      valid[39] = 1;
      outs[39] = outs[38];
    end
    else begin
      if (decode_signal[38]) begin
        valid[39] = 1;
        outs[39] = 38;
      end
      else begin
        valid[39] = 0;
        outs[39] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[39]) begin
      valid[40] = 1;
      outs[40] = outs[39];
    end
    else begin
      if (decode_signal[39]) begin
        valid[40] = 1;
        outs[40] = 39;
      end
      else begin
        valid[40] = 0;
        outs[40] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[40]) begin
      valid[41] = 1;
      outs[41] = outs[40];
    end
    else begin
      if (decode_signal[40]) begin
        valid[41] = 1;
        outs[41] = 40;
      end
      else begin
        valid[41] = 0;
        outs[41] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[41]) begin
      valid[42] = 1;
      outs[42] = outs[41];
    end
    else begin
      if (decode_signal[41]) begin
        valid[42] = 1;
        outs[42] = 41;
      end
      else begin
        valid[42] = 0;
        outs[42] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[42]) begin
      valid[43] = 1;
      outs[43] = outs[42];
    end
    else begin
      if (decode_signal[42]) begin
        valid[43] = 1;
        outs[43] = 42;
      end
      else begin
        valid[43] = 0;
        outs[43] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[43]) begin
      valid[44] = 1;
      outs[44] = outs[43];
    end
    else begin
      if (decode_signal[43]) begin
        valid[44] = 1;
        outs[44] = 43;
      end
      else begin
        valid[44] = 0;
        outs[44] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[44]) begin
      valid[45] = 1;
      outs[45] = outs[44];
    end
    else begin
      if (decode_signal[44]) begin
        valid[45] = 1;
        outs[45] = 44;
      end
      else begin
        valid[45] = 0;
        outs[45] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[45]) begin
      valid[46] = 1;
      outs[46] = outs[45];
    end
    else begin
      if (decode_signal[45]) begin
        valid[46] = 1;
        outs[46] = 45;
      end
      else begin
        valid[46] = 0;
        outs[46] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[46]) begin
      valid[47] = 1;
      outs[47] = outs[46];
    end
    else begin
      if (decode_signal[46]) begin
        valid[47] = 1;
        outs[47] = 46;
      end
      else begin
        valid[47] = 0;
        outs[47] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[47]) begin
      valid[48] = 1;
      outs[48] = outs[47];
    end
    else begin
      if (decode_signal[47]) begin
        valid[48] = 1;
        outs[48] = 47;
      end
      else begin
        valid[48] = 0;
        outs[48] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[48]) begin
      valid[49] = 1;
      outs[49] = outs[48];
    end
    else begin
      if (decode_signal[48]) begin
        valid[49] = 1;
        outs[49] = 48;
      end
      else begin
        valid[49] = 0;
        outs[49] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[49]) begin
      valid[50] = 1;
      outs[50] = outs[49];
    end
    else begin
      if (decode_signal[49]) begin
        valid[50] = 1;
        outs[50] = 49;
      end
      else begin
        valid[50] = 0;
        outs[50] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[50]) begin
      valid[51] = 1;
      outs[51] = outs[50];
    end
    else begin
      if (decode_signal[50]) begin
        valid[51] = 1;
        outs[51] = 50;
      end
      else begin
        valid[51] = 0;
        outs[51] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[51]) begin
      valid[52] = 1;
      outs[52] = outs[51];
    end
    else begin
      if (decode_signal[51]) begin
        valid[52] = 1;
        outs[52] = 51;
      end
      else begin
        valid[52] = 0;
        outs[52] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[52]) begin
      valid[53] = 1;
      outs[53] = outs[52];
    end
    else begin
      if (decode_signal[52]) begin
        valid[53] = 1;
        outs[53] = 52;
      end
      else begin
        valid[53] = 0;
        outs[53] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[53]) begin
      valid[54] = 1;
      outs[54] = outs[53];
    end
    else begin
      if (decode_signal[53]) begin
        valid[54] = 1;
        outs[54] = 53;
      end
      else begin
        valid[54] = 0;
        outs[54] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[54]) begin
      valid[55] = 1;
      outs[55] = outs[54];
    end
    else begin
      if (decode_signal[54]) begin
        valid[55] = 1;
        outs[55] = 54;
      end
      else begin
        valid[55] = 0;
        outs[55] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[55]) begin
      valid[56] = 1;
      outs[56] = outs[55];
    end
    else begin
      if (decode_signal[55]) begin
        valid[56] = 1;
        outs[56] = 55;
      end
      else begin
        valid[56] = 0;
        outs[56] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[56]) begin
      valid[57] = 1;
      outs[57] = outs[56];
    end
    else begin
      if (decode_signal[56]) begin
        valid[57] = 1;
        outs[57] = 56;
      end
      else begin
        valid[57] = 0;
        outs[57] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[57]) begin
      valid[58] = 1;
      outs[58] = outs[57];
    end
    else begin
      if (decode_signal[57]) begin
        valid[58] = 1;
        outs[58] = 57;
      end
      else begin
        valid[58] = 0;
        outs[58] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[58]) begin
      valid[59] = 1;
      outs[59] = outs[58];
    end
    else begin
      if (decode_signal[58]) begin
        valid[59] = 1;
        outs[59] = 58;
      end
      else begin
        valid[59] = 0;
        outs[59] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[59]) begin
      valid[60] = 1;
      outs[60] = outs[59];
    end
    else begin
      if (decode_signal[59]) begin
        valid[60] = 1;
        outs[60] = 59;
      end
      else begin
        valid[60] = 0;
        outs[60] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[60]) begin
      valid[61] = 1;
      outs[61] = outs[60];
    end
    else begin
      if (decode_signal[60]) begin
        valid[61] = 1;
        outs[61] = 60;
      end
      else begin
        valid[61] = 0;
        outs[61] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[61]) begin
      valid[62] = 1;
      outs[62] = outs[61];
    end
    else begin
      if (decode_signal[61]) begin
        valid[62] = 1;
        outs[62] = 61;
      end
      else begin
        valid[62] = 0;
        outs[62] = 0;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_decode(n=i + 1, i=i):
  //         if s.valid[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = s.outs[i]
  //         elif s.decode_signal[i]:
  //           s.valid[n].v = 1
  //           s.outs[n].v = i
  //         else:
  //           s.valid[n].v = 0
  //           s.outs[n].v = 0

  // logic for handle_decode()
  always @ (*) begin
    if (valid[62]) begin
      valid[63] = 1;
      outs[63] = outs[62];
    end
    else begin
      if (decode_signal[62]) begin
        valid[63] = 1;
        outs[63] = 62;
      end
      else begin
        valid[63] = 0;
        outs[63] = 0;
      end
    end
  end


endmodule // PriorityDecoder_0x2e5c0266b41857fd

//-----------------------------------------------------------------------------
// KillNotifier_0x40986fce6fe74c56
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.kill_unit {"KillArgType": 5}
// PyMTL: verilator_xinit = zeros
module KillNotifier_0x40986fce6fe74c56
(
  input  logic [   4:0] check_kill_kill,
  input  logic [   0:0] clk,
  output logic [   4:0] kill_notify_msg,
  input  logic [   0:0] reset
);

  // signal connections
  assign kill_notify_msg = check_kill_kill;



endmodule // KillNotifier_0x40986fce6fe74c56

//-----------------------------------------------------------------------------
// PipelineArbiter_0x311a0425acf3e6db
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.pipeline_arbiter {"clients": ["alu", "csr", "branch"], "interface": "peek <R> () -> (msg: Bits(146)); take <C> () -> ()"}
// PyMTL: verilator_xinit = zeros
module PipelineArbiter_0x311a0425acf3e6db
(
  input  logic [ 145:0] alu_peek_msg,
  input  logic [   0:0] alu_peek_rdy,
  output logic [   0:0] alu_take_call,
  input  logic [ 145:0] branch_peek_msg,
  input  logic [   0:0] branch_peek_rdy,
  output logic [   0:0] branch_take_call,
  input  logic [   0:0] clk,
  input  logic [ 145:0] csr_peek_msg,
  input  logic [   0:0] csr_peek_rdy,
  output logic [   0:0] csr_take_call,
  output logic [ 145:0] peek_msg,
  output logic  [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // logic declarations
  logic   [ 145:0] index_peek_msg$000;
  logic   [ 145:0] index_peek_msg$001;
  logic   [ 145:0] index_peek_msg$002;
  logic   [   0:0] index_take_call$000;
  logic   [   0:0] index_take_call$001;
  logic   [   0:0] index_take_call$002;
  logic   [   0:0] index_peek_rdy$000;
  logic   [   0:0] index_peek_rdy$001;
  logic   [   0:0] index_peek_rdy$002;


  // arb temporaries
  logic   [   2:0] arb$grant_reqs;
  logic   [   0:0] arb$clk;
  logic   [   0:0] arb$reset;
  logic   [   2:0] arb$grant_grant;

  RoundRobinArbiter_0x5f763cfe8f4295d1 arb
  (
    .grant_reqs  ( arb$grant_reqs ),
    .clk         ( arb$clk ),
    .reset       ( arb$reset ),
    .grant_grant ( arb$grant_grant )
  );

  // mux temporaries
  logic   [ 145:0] mux$mux_default;
  logic   [ 145:0] mux$mux_in_$000;
  logic   [ 145:0] mux$mux_in_$001;
  logic   [ 145:0] mux$mux_in_$002;
  logic   [   0:0] mux$clk;
  logic   [   0:0] mux$reset;
  logic   [   2:0] mux$mux_select;
  logic   [ 145:0] mux$mux_out;
  logic   [   0:0] mux$mux_matched;

  CaseMux_0x2a6155b79f50b353 mux
  (
    .mux_default ( mux$mux_default ),
    .mux_in_$000 ( mux$mux_in_$000 ),
    .mux_in_$001 ( mux$mux_in_$001 ),
    .mux_in_$002 ( mux$mux_in_$002 ),
    .clk         ( mux$clk ),
    .reset       ( mux$reset ),
    .mux_select  ( mux$mux_select ),
    .mux_out     ( mux$mux_out ),
    .mux_matched ( mux$mux_matched )
  );

  // signal connections
  assign alu_take_call      = index_take_call$000;
  assign arb$clk            = clk;
  assign arb$grant_reqs[0]  = index_peek_rdy$000;
  assign arb$grant_reqs[1]  = index_peek_rdy$001;
  assign arb$grant_reqs[2]  = index_peek_rdy$002;
  assign arb$reset          = reset;
  assign branch_take_call   = index_take_call$002;
  assign csr_take_call      = index_take_call$001;
  assign index_peek_msg$000 = alu_peek_msg;
  assign index_peek_msg$001 = csr_peek_msg;
  assign index_peek_msg$002 = branch_peek_msg;
  assign index_peek_rdy$000 = alu_peek_rdy;
  assign index_peek_rdy$001 = csr_peek_rdy;
  assign index_peek_rdy$002 = branch_peek_rdy;
  assign mux$clk            = clk;
  assign mux$mux_default    = 146'd0;
  assign mux$mux_in_$000    = index_peek_msg$000;
  assign mux$mux_in_$001    = index_peek_msg$001;
  assign mux$mux_in_$002    = index_peek_msg$002;
  assign mux$mux_select     = arb$grant_grant;
  assign mux$reset          = reset;
  assign peek_msg           = mux$mux_out;

  // array declarations
  logic    [   0:0] index_take_call[0:2];
  assign index_take_call$000 = index_take_call[  0];
  assign index_take_call$001 = index_take_call[  1];
  assign index_take_call$002 = index_take_call[  2];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_ready():
  //       s.peek_rdy.v = (s.arb.grant_grant != 0)

  // logic for compute_ready()
  always @ (*) begin
    peek_rdy = (arb$grant_grant != 0);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_call(i=i):
  //         s.index_take_call[i].v = s.arb.grant_grant[i] & s.take_call

  // logic for compute_call()
  always @ (*) begin
    index_take_call[0] = (arb$grant_grant[0]&take_call);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_call(i=i):
  //         s.index_take_call[i].v = s.arb.grant_grant[i] & s.take_call

  // logic for compute_call()
  always @ (*) begin
    index_take_call[1] = (arb$grant_grant[1]&take_call);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute_call(i=i):
  //         s.index_take_call[i].v = s.arb.grant_grant[i] & s.take_call

  // logic for compute_call()
  always @ (*) begin
    index_take_call[2] = (arb$grant_grant[2]&take_call);
  end


endmodule // PipelineArbiter_0x311a0425acf3e6db

//-----------------------------------------------------------------------------
// RoundRobinArbiter_0x5f763cfe8f4295d1
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.arbiters {"interface": "grant (reqs: Bits(3)) -> (grant: Bits(3))"}
// PyMTL: verilator_xinit = zeros
module RoundRobinArbiter_0x5f763cfe8f4295d1
(
  input  logic [   0:0] clk,
  output logic [   2:0] grant_grant,
  input  logic [   2:0] grant_reqs,
  input  logic [   0:0] reset
);

  // register declarations
  logic    [   2:0] final_grant;
  logic    [   2:0] masked_arb$grant_reqs;

  // masker temporaries
  logic   [   0:0] masker$clk;
  logic   [   0:0] masker$reset;
  logic   [   2:0] masker$mask_in_;
  logic   [   2:0] masker$mask_out;

  ThermometerMask_0x4e5c8d2b7524bd9b masker
  (
    .clk      ( masker$clk ),
    .reset    ( masker$reset ),
    .mask_in_ ( masker$mask_in_ ),
    .mask_out ( masker$mask_out )
  );

  // raw_arb temporaries
  logic   [   2:0] raw_arb$grant_reqs;
  logic   [   0:0] raw_arb$clk;
  logic   [   0:0] raw_arb$reset;
  logic   [   2:0] raw_arb$grant_grant;

  PriorityArbiter_0x5f763cfe8f4295d1 raw_arb
  (
    .grant_reqs  ( raw_arb$grant_reqs ),
    .clk         ( raw_arb$clk ),
    .reset       ( raw_arb$reset ),
    .grant_grant ( raw_arb$grant_grant )
  );

  // masked_arb temporaries
  logic   [   0:0] masked_arb$clk;
  logic   [   0:0] masked_arb$reset;
  logic   [   2:0] masked_arb$grant_grant;

  PriorityArbiter_0x5f763cfe8f4295d1 masked_arb
  (
    .grant_reqs  ( masked_arb$grant_reqs ),
    .clk         ( masked_arb$clk ),
    .reset       ( masked_arb$reset ),
    .grant_grant ( masked_arb$grant_grant )
  );

  // mask temporaries
  logic   [   0:0] mask$clk;
  logic   [   2:0] mask$write_data;
  logic   [   0:0] mask$reset;
  logic   [   2:0] mask$read_data;

  Register_0x3e6a7278e29c371 mask
  (
    .clk        ( mask$clk ),
    .write_data ( mask$write_data ),
    .reset      ( mask$reset ),
    .read_data  ( mask$read_data )
  );

  // signal connections
  assign grant_grant        = final_grant;
  assign mask$clk           = clk;
  assign mask$reset         = reset;
  assign mask$write_data    = final_grant;
  assign masked_arb$clk     = clk;
  assign masked_arb$reset   = reset;
  assign masker$clk         = clk;
  assign masker$mask_in_    = mask$read_data;
  assign masker$reset       = reset;
  assign raw_arb$clk        = clk;
  assign raw_arb$grant_reqs = grant_reqs;
  assign raw_arb$reset      = reset;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute():
  //       s.masked_arb.grant_reqs.v = s.grant_reqs & s.masker.mask_out
  //       if s.masked_arb.grant_grant == 0:
  //         s.final_grant.v = s.raw_arb.grant_grant
  //       else:
  //         s.final_grant.v = s.masked_arb.grant_grant

  // logic for compute()
  always @ (*) begin
    masked_arb$grant_reqs = (grant_reqs&masker$mask_out);
    if ((masked_arb$grant_grant == 0)) begin
      final_grant = raw_arb$grant_grant;
    end
    else begin
      final_grant = masked_arb$grant_grant;
    end
  end


endmodule // RoundRobinArbiter_0x5f763cfe8f4295d1

//-----------------------------------------------------------------------------
// ThermometerMask_0x4e5c8d2b7524bd9b
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.thermometer_mask {"interface": "mask (in_: Bits(3)) -> (out: Bits(3))"}
// PyMTL: verilator_xinit = zeros
module ThermometerMask_0x4e5c8d2b7524bd9b
(
  input  logic [   0:0] clk,
  input  logic [   2:0] mask_in_,
  output logic  [   2:0] mask_out,
  input  logic [   0:0] reset
);



  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute():
  //       s.mask_out.v = s.mask_in_ ^ (s.mask_in_ - 1)
  //       s.mask_out.v = s.mask_out if s.mask_in_ == 0 else ~s.mask_out
  //       s.mask_out.v = s.mask_out | s.mask_in_

  // logic for compute()
  always @ (*) begin
    mask_out = (mask_in_^(mask_in_-1));
    mask_out = (mask_in_ == 0) ? mask_out : ~mask_out;
    mask_out = (mask_out|mask_in_);
  end


endmodule // ThermometerMask_0x4e5c8d2b7524bd9b

//-----------------------------------------------------------------------------
// PriorityArbiter_0x5f763cfe8f4295d1
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.arbiters {"interface": "grant (reqs: Bits(3)) -> (grant: Bits(3))"}
// PyMTL: verilator_xinit = zeros
module PriorityArbiter_0x5f763cfe8f4295d1
(
  input  logic [   0:0] clk,
  output logic  [   2:0] grant_grant,
  input  logic [   2:0] grant_reqs,
  input  logic [   0:0] reset
);



  // PYMTL SOURCE:
  //
  // @s.combinational
  // def compute():
  //       # PYMTL_BROKEN unary - translates but does not simulate
  //       s.grant_grant.v = s.grant_reqs & (0 - s.grant_reqs)

  // logic for compute()
  always @ (*) begin
    grant_grant = (grant_reqs&(0-grant_reqs));
  end


endmodule // PriorityArbiter_0x5f763cfe8f4295d1

//-----------------------------------------------------------------------------
// Register_0x3e6a7278e29c371
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(3)); write (data: Bits(3)) -> ()", "reset_value": 0}
// PyMTL: verilator_xinit = zeros
module Register_0x3e6a7278e29c371
(
  input  logic [   0:0] clk,
  output logic [   2:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   2:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [   2:0] reg_value;

  // localparam declarations
  localparam reset_value = 0;

  // signal connections
  assign read_data = reg_value;
  assign update    = 1'd1;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.reset:
  //           s.reg_value.n = reset_value
  //         elif s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      reg_value <= reset_value;
    end
    else begin
      if (update) begin
        reg_value <= write_data;
      end
      else begin
      end
    end
  end


endmodule // Register_0x3e6a7278e29c371

//-----------------------------------------------------------------------------
// CaseMux_0x2a6155b79f50b353
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.case_mux {"interface": "mux (default: Bits(146), in_: Bits(146) [3], select: Bits(3)) -> (out: Bits(146), matched: Bits(1))", "svalues": [1, 2, 4]}
// PyMTL: verilator_xinit = zeros
module CaseMux_0x2a6155b79f50b353
(
  input  logic [   0:0] clk,
  input  logic [ 145:0] mux_default,
  input  logic [ 145:0] mux_in_$000,
  input  logic [ 145:0] mux_in_$001,
  input  logic [ 145:0] mux_in_$002,
  output logic [   0:0] mux_matched,
  output logic [ 145:0] mux_out,
  input  logic [   2:0] mux_select,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [ 145:0] out_chain$000;
  logic   [ 145:0] out_chain$001;
  logic   [ 145:0] out_chain$002;
  logic   [ 145:0] out_chain$003;
  logic   [   0:0] valid_chain$000;
  logic   [   0:0] valid_chain$001;
  logic   [   0:0] valid_chain$002;
  logic   [   0:0] valid_chain$003;


  // signal connections
  assign mux_matched     = valid_chain$003;
  assign mux_out         = out_chain$003;
  assign valid_chain$000 = 1'd0;

  // array declarations
  logic   [ 145:0] mux_in_[0:2];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  logic    [ 145:0] out_chain[0:3];
  assign out_chain$000 = out_chain[  0];
  assign out_chain$001 = out_chain[  1];
  assign out_chain$002 = out_chain[  2];
  assign out_chain$003 = out_chain[  3];
  logic    [   0:0] valid_chain[0:3];
  assign valid_chain$000 = valid_chain[  0];
  assign valid_chain$001 = valid_chain[  1];
  assign valid_chain$002 = valid_chain[  2];
  assign valid_chain$003 = valid_chain[  3];

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def connect_is_broken():
  //       s.out_chain[0].v = s.mux_default

  // logic for connect_is_broken()
  always @ (*) begin
    out_chain[0] = mux_default;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 1)) begin
      out_chain[1] = mux_in_[0];
      valid_chain[1] = 1;
    end
    else begin
      out_chain[1] = out_chain[0];
      valid_chain[1] = valid_chain[0];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 2)) begin
      out_chain[2] = mux_in_[1];
      valid_chain[2] = 1;
    end
    else begin
      out_chain[2] = out_chain[1];
      valid_chain[2] = valid_chain[1];
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def chain(curr=i + 1, last=i, svalue=int(svalue)):
  //         if s.mux_select == svalue:
  //           s.out_chain[curr].v = s.mux_in_[last]
  //           s.valid_chain[curr].v = 1
  //         else:
  //           s.out_chain[curr].v = s.out_chain[last]
  //           s.valid_chain[curr].v = s.valid_chain[last]

  // logic for chain()
  always @ (*) begin
    if ((mux_select == 4)) begin
      out_chain[3] = mux_in_[2];
      valid_chain[3] = 1;
    end
    else begin
      out_chain[3] = out_chain[2];
      valid_chain[3] = valid_chain[2];
    end
  end


endmodule // CaseMux_0x2a6155b79f50b353

//-----------------------------------------------------------------------------
// ControlFlowManager_0x734ebf4161405225
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.controlflow {"cflow_interface": "check_kill () -> (kill: Bits(5)); check_redirect () -> (redirect: Bits(1), target: Bits(64)); commit <C> (status: Bits(2)) -> (); get_head <R> () -> (seq: Bits(4)); redirect <C> (spec_idx: Bits(1), force: Bits(1), target: Bits(64), seq: Bits(4)) -> (); register <C> (pc: Bits(64), speculative: Bits(1), serialize: Bits(1), pc_succ: Bits(64)) -> (branch_mask: Bits(2), spec_idx: Bits(1), seq: Bits(4), success: Bits(1))", "reset_vector": 64, "trap_vector": 0}
// PyMTL: verilator_xinit = zeros
module ControlFlowManager_0x734ebf4161405225
(
  output logic [   4:0] check_kill_kill,
  output logic  [   0:0] check_redirect_redirect,
  output logic  [  63:0] check_redirect_target,
  input  logic [   0:0] clk,
  input  logic [   0:0] commit_call,
  input  logic [   1:0] commit_status,
  output logic  [   0:0] dflow_free_snapshot_call,
  output logic [   0:0] dflow_free_snapshot_id_,
  output logic [   0:0] dflow_restore_call,
  output logic [   0:0] dflow_restore_source_id,
  output logic  [   0:0] dflow_rollback_call,
  output logic [   0:0] dflow_snapshot_call,
  input  logic [   0:0] dflow_snapshot_id_,
  input  logic [   0:0] dflow_snapshot_rdy,
  output logic  [   0:0] get_head_rdy,
  output logic [   3:0] get_head_seq,
  input  logic [   0:0] redirect_call,
  input  logic [   0:0] redirect_force,
  input  logic [   3:0] redirect_seq,
  input  logic [   0:0] redirect_spec_idx,
  input  logic [  63:0] redirect_target,
  output logic [   1:0] register_branch_mask,
  input  logic [   0:0] register_call,
  input  logic [  63:0] register_pc,
  input  logic [  63:0] register_pc_succ,
  output logic [   3:0] register_seq,
  input  logic [   0:0] register_serialize,
  output logic [   0:0] register_spec_idx,
  input  logic [   0:0] register_speculative,
  output logic [   0:0] register_success,
  input  logic [   0:0] reset
);

  // register declarations
  logic    [   0:0] bmask$write_call;
  logic    [   1:0] bmask_curr_;
  logic    [   1:0] bmask_next_;
  logic    [   1:0] clear_mask_;
  logic    [   0:0] commit_redirect_;
  logic    [  63:0] commit_redirect_target_;
  logic    [   0:0] empty_;
  logic    [   0:0] full_;
  logic    [   0:0] head$write_call;
  logic    [   3:0] head$write_data;
  logic    [   3:0] head_next;
  logic    [   3:0] head_tail_delta;
  logic    [   1:0] kill_mask_;
  logic    [   0:0] num$write_call;
  logic    [   4:0] num$write_data;
  logic    [   0:0] redirect_;
  logic    [  63:0] redirect_target_;
  logic    [   0:0] register_success_;
  logic    [   0:0] reset_redirect_valid_;
  logic    [   0:0] serial$write_call;
  logic    [   0:0] serial$write_data;
  logic    [   0:0] spec_register_success_;
  logic    [   0:0] tail$write_call;
  logic    [   3:0] tail$write_data;

  // localparam declarations
  localparam PIPELINE_MSG_STATUS_VALID = 2'd0;
  localparam max_entries = 16;
  localparam reset_vector = 64'd512;
  localparam trap_vector = 0;

  // tail temporaries
  logic   [   0:0] tail$clk;
  logic   [   0:0] tail$reset;
  logic   [   3:0] tail$read_data;

  Register_0x5d4baebedb8e9d8 tail
  (
    .clk        ( tail$clk ),
    .write_call ( tail$write_call ),
    .write_data ( tail$write_data ),
    .reset      ( tail$reset ),
    .read_data  ( tail$read_data )
  );

  // bmask_alloc temporaries
  logic   [   0:0] bmask_alloc$encode_call;
  logic   [   0:0] bmask_alloc$clk;
  logic   [   0:0] bmask_alloc$reset;
  logic   [   0:0] bmask_alloc$encode_number;
  logic   [   1:0] bmask_alloc$encode_onehot;

  OneHotEncoder_0x6ddac805079c9f17 bmask_alloc
  (
    .encode_call   ( bmask_alloc$encode_call ),
    .clk           ( bmask_alloc$clk ),
    .reset         ( bmask_alloc$reset ),
    .encode_number ( bmask_alloc$encode_number ),
    .encode_onehot ( bmask_alloc$encode_onehot )
  );

  // redirect_mask temporaries
  logic   [   0:0] redirect_mask$clk;
  logic   [   0:0] redirect_mask$reset;
  logic   [   0:0] redirect_mask$encode_number;
  logic   [   1:0] redirect_mask$encode_onehot;

  OneHotEncoder_0x62af1c1ff9e32b51 redirect_mask
  (
    .clk           ( redirect_mask$clk ),
    .reset         ( redirect_mask$reset ),
    .encode_number ( redirect_mask$encode_number ),
    .encode_onehot ( redirect_mask$encode_onehot )
  );

  // num temporaries
  logic   [   0:0] num$clk;
  logic   [   0:0] num$reset;
  logic   [   4:0] num$read_data;

  Register_0xae4a367f21f784a num
  (
    .clk        ( num$clk ),
    .write_call ( num$write_call ),
    .write_data ( num$write_data ),
    .reset      ( num$reset ),
    .read_data  ( num$read_data )
  );

  // head temporaries
  logic   [   0:0] head$clk;
  logic   [   0:0] head$reset;
  logic   [   3:0] head$read_data;

  Register_0x5d4baebedb8e9d8 head
  (
    .clk        ( head$clk ),
    .write_call ( head$write_call ),
    .write_data ( head$write_data ),
    .reset      ( head$reset ),
    .read_data  ( head$read_data )
  );

  // pc_pred temporaries
  logic   [   0:0] pc_pred$clk;
  logic   [   0:0] pc_pred$write_addr$000;
  logic   [   0:0] pc_pred$read_addr$000;
  logic   [   0:0] pc_pred$write_call$000;
  logic   [  63:0] pc_pred$write_data$000;
  logic   [   0:0] pc_pred$reset;
  logic   [  63:0] pc_pred$read_data$000;

  AsynchronousRAM_0x7bb0942938a43a9 pc_pred
  (
    .clk            ( pc_pred$clk ),
    .write_addr$000 ( pc_pred$write_addr$000 ),
    .read_addr$000  ( pc_pred$read_addr$000 ),
    .write_call$000 ( pc_pred$write_call$000 ),
    .write_data$000 ( pc_pred$write_data$000 ),
    .reset          ( pc_pred$reset ),
    .read_data$000  ( pc_pred$read_data$000 )
  );

  // serial temporaries
  logic   [   0:0] serial$clk;
  logic   [   0:0] serial$reset;
  logic   [   0:0] serial$read_data;

  Register_0x19ffe7c045ca5b3a serial
  (
    .clk        ( serial$clk ),
    .write_call ( serial$write_call ),
    .write_data ( serial$write_data ),
    .reset      ( serial$reset ),
    .read_data  ( serial$read_data )
  );

  // bmask temporaries
  logic   [   0:0] bmask$clk;
  logic   [   1:0] bmask$write_data;
  logic   [   0:0] bmask$reset;
  logic   [   1:0] bmask$read_data;

  Register_0x60b9ec19bb3fa768 bmask
  (
    .clk        ( bmask$clk ),
    .write_call ( bmask$write_call ),
    .write_data ( bmask$write_data ),
    .reset      ( bmask$reset ),
    .read_data  ( bmask$read_data )
  );

  // signal connections
  assign bmask$clk                   = clk;
  assign bmask$reset                 = reset;
  assign bmask$write_data            = bmask_next_;
  assign bmask_alloc$clk             = clk;
  assign bmask_alloc$encode_call     = spec_register_success_;
  assign bmask_alloc$encode_number   = dflow_snapshot_id_;
  assign bmask_alloc$reset           = reset;
  assign check_kill_kill[0:0]        = redirect_force;
  assign check_kill_kill[2:1]        = kill_mask_;
  assign check_kill_kill[4:3]        = clear_mask_;
  assign dflow_free_snapshot_id_     = redirect_spec_idx;
  assign dflow_restore_call          = redirect_;
  assign dflow_restore_source_id     = redirect_spec_idx;
  assign dflow_snapshot_call         = spec_register_success_;
  assign get_head_seq                = head$read_data;
  assign head$clk                    = clk;
  assign head$reset                  = reset;
  assign num$clk                     = clk;
  assign num$reset                   = reset;
  assign pc_pred$clk                 = clk;
  assign pc_pred$read_addr$000       = redirect_spec_idx;
  assign pc_pred$reset               = reset;
  assign pc_pred$write_addr$000      = dflow_snapshot_id_;
  assign pc_pred$write_call$000      = spec_register_success_;
  assign pc_pred$write_data$000      = register_pc_succ;
  assign redirect_mask$clk           = clk;
  assign redirect_mask$encode_number = redirect_spec_idx;
  assign redirect_mask$reset         = reset;
  assign register_branch_mask        = bmask_curr_;
  assign register_seq                = tail$read_data;
  assign register_spec_idx           = dflow_snapshot_id_;
  assign register_success            = register_success_;
  assign serial$clk                  = clk;
  assign serial$reset                = reset;
  assign tail$clk                    = clk;
  assign tail$reset                  = reset;

  // array declarations
  logic   [  63:0] pc_pred$read_data[0:0];
  assign pc_pred$read_data[  0] = pc_pred$read_data$000;

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def handle_reset():
  //       s.reset_redirect_valid_.n = s.reset

  // logic for handle_reset()
  always @ (posedge clk) begin
    reset_redirect_valid_ <= reset;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def prioritry_redirect():
  //       s.check_redirect_redirect.v = s.reset_redirect_valid_ or s.commit_redirect_ or s.redirect_
  //       s.check_redirect_target.v = 0
  //       if s.reset_redirect_valid_:
  //         s.check_redirect_target.v = reset_vector
  //       elif s.commit_redirect_:
  //         s.check_redirect_target.v = s.commit_redirect_target_
  //       else:  # s.redirect_
  //         s.check_redirect_target.v = s.redirect_target_

  // logic for prioritry_redirect()
  always @ (*) begin
    check_redirect_redirect = (reset_redirect_valid_||commit_redirect_||redirect_);
    check_redirect_target = 0;
    if (reset_redirect_valid_) begin
      check_redirect_target = reset_vector;
    end
    else begin
      if (commit_redirect_) begin
        check_redirect_target = commit_redirect_target_;
      end
      else begin
        check_redirect_target = redirect_target_;
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_serial():
  //       s.serial.write_call.v = ((s.register_success and s.register_serialize) or
  //                                (s.serial.read_data and s.commit_call))
  //       s.serial.write_data.v = not s.serial.read_data  #  we are always inverting it

  // logic for set_serial()
  always @ (*) begin
    serial$write_call = ((register_success&&register_serialize)||(serial$read_data&&commit_call));
    serial$write_data = !serial$read_data;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_redirection():
  //       # These are set after a redirect call
  //       s.kill_mask_.v = 0
  //       s.clear_mask_.v = 0
  //       s.redirect_.v = 0
  //       s.redirect_target_.v = 0
  //       s.dflow_free_snapshot_call.v = 0
  //       if s.redirect_call:
  //         # Free the snapshot
  //         s.dflow_free_snapshot_call.v = 1
  //         # Look up if the predicted PC saved during register is correct
  //         s.redirect_.v = s.redirect_target != s.pc_pred.read_data[
  //             0] or s.redirect_force
  //         if s.redirect_:
  //           s.kill_mask_.v = s.redirect_mask.encode_onehot
  //           s.redirect_target_.v = s.redirect_target
  //         else:
  //           s.clear_mask_.v = s.redirect_mask.encode_onehot

  // logic for handle_redirection()
  always @ (*) begin
    kill_mask_ = 0;
    clear_mask_ = 0;
    redirect_ = 0;
    redirect_target_ = 0;
    dflow_free_snapshot_call = 0;
    if (redirect_call) begin
      dflow_free_snapshot_call = 1;
      redirect_ = ((redirect_target != pc_pred$read_data[0])||redirect_force);
      if (redirect_) begin
        kill_mask_ = redirect_mask$encode_onehot;
        redirect_target_ = redirect_target;
      end
      else begin
        clear_mask_ = redirect_mask$encode_onehot;
      end
    end
    else begin
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_bmask():
  //       s.bmask.write_call.v = s.spec_register_success_ or s.redirect_call or s.commit_redirect_
  //       # Update the current branch mask
  //       s.bmask_curr_.v = s.bmask.read_data.v & (~(s.kill_mask_ | s.clear_mask_))
  //       s.bmask_next_.v = s.bmask_curr_
  //       if s.commit_redirect_:
  //         s.bmask_next_.v = 0
  //       elif s.register_speculative:
  //         s.bmask_next_.v = s.bmask_curr_ | s.bmask_alloc.encode_onehot

  // logic for handle_bmask()
  always @ (*) begin
    bmask$write_call = (spec_register_success_||redirect_call||commit_redirect_);
    bmask_curr_ = (bmask$read_data&~(kill_mask_|clear_mask_));
    bmask_next_ = bmask_curr_;
    if (commit_redirect_) begin
      bmask_next_ = 0;
    end
    else begin
      if (register_speculative) begin
        bmask_next_ = (bmask_curr_|bmask_alloc$encode_onehot);
      end
      else begin
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_register():
  //       # TODO handle speculative
  //       s.register_success_.v = 0
  //       s.spec_register_success_.v = 0
  //       if s.register_call:
  //         s.register_success_.v = (not s.full_ and (not s.register_speculative or
  //                                                   s.dflow_snapshot_rdy) and
  //                                  (not s.register_serialize or s.empty_) and
  //                                  not s.serial.read_data)
  //
  //         s.spec_register_success_.v = s.register_success_.v and s.register_speculative

  // logic for handle_register()
  always @ (*) begin
    register_success_ = 0;
    spec_register_success_ = 0;
    if (register_call) begin
      register_success_ = (!full_&&(!register_speculative||dflow_snapshot_rdy)&&(!register_serialize||empty_)&&!serial$read_data);
      spec_register_success_ = (register_success_&&register_speculative);
    end
    else begin
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_commit():
  //       s.dflow_rollback_call.v = 0
  //       #s.dflow_free_snapshot_call.v = 0
  //       s.commit_redirect_.v = 0
  //       s.commit_redirect_target_.v = 0
  //       # If we are committing there are a couple cases
  //       if s.commit_call:
  //         # Jump to exception handler
  //         if s.commit_status != PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID:
  //           # TODO jump to proper handler
  //           s.commit_redirect_target_.v = trap_vector
  //           s.commit_redirect_.v = 1
  //           s.dflow_rollback_call.v = 1

  // logic for handle_commit()
  always @ (*) begin
    dflow_rollback_call = 0;
    commit_redirect_ = 0;
    commit_redirect_target_ = 0;
    if (commit_call) begin
      if ((commit_status != PIPELINE_MSG_STATUS_VALID)) begin
        commit_redirect_target_ = trap_vector;
        commit_redirect_ = 1;
        dflow_rollback_call = 1;
      end
      else begin
      end
    end
    else begin
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_get_head_rdy():
  //       s.get_head_rdy.v = not s.empty_

  // logic for set_get_head_rdy()
  always @ (*) begin
    get_head_rdy = !empty_;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_flags():
  //       s.full_.v = s.num.read_data == max_entries
  //       s.empty_.v = s.num.read_data == 0

  // logic for set_flags()
  always @ (*) begin
    full_ = (num$read_data == max_entries);
    empty_ = (num$read_data == 0);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_tail():
  //       s.tail.write_call.v = s.register_success or s.commit_redirect_ or s.redirect_
  //       if s.commit_redirect_:
  //         # On an exception, the tail = head + 1, since head will be incremented
  //         s.tail.write_data.v = s.head.read_data + 1
  //       elif s.redirect_:
  //         s.tail.write_data.v = s.redirect_seq + 1  # Note: Tail is exclusive
  //       else:
  //         s.tail.write_data.v = s.tail.read_data + 1

  // logic for update_tail()
  always @ (*) begin
    tail$write_call = (register_success||commit_redirect_||redirect_);
    if (commit_redirect_) begin
      tail$write_data = (head$read_data+1);
    end
    else begin
      if (redirect_) begin
        tail$write_data = (redirect_seq+1);
      end
      else begin
        tail$write_data = (tail$read_data+1);
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_head():
  //       s.head_next.v = s.head.read_data + 1 if s.commit_call else s.head.read_data
  //       s.head.write_call.v = s.commit_call
  //       s.head.write_data.v = s.head_next

  // logic for update_head()
  always @ (*) begin
    head_next = commit_call ? (head$read_data+1) : head$read_data;
    head$write_call = commit_call;
    head$write_data = head_next;
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def update_num(seqp1=seqidx_nbits + 1):
  //       s.head_tail_delta.v = s.tail.write_data - s.head_next
  //       s.num.write_call.v = s.tail.write_call or s.head.write_call
  //       s.num.write_data.v = s.num.read_data
  //       if s.commit_redirect_:
  //         s.num.write_data.v = 0  # An exception clears everything
  //       elif s.redirect_:
  //         s.num.write_data.v = max_entries if s.head_tail_delta == 0 else zext(
  //             s.head_tail_delta, seqp1)
  //       elif s.register_success ^ s.commit_call:
  //         if s.register_success:
  //           s.num.write_data.v = s.num.read_data + 1
  //         elif s.commit_call:
  //           s.num.write_data.v = s.num.read_data - 1

  // logic for update_num()
  always @ (*) begin
    head_tail_delta = (tail$write_data-head_next);
    num$write_call = (tail$write_call||head$write_call);
    num$write_data = num$read_data;
    if (commit_redirect_) begin
      num$write_data = 0;
    end
    else begin
      if (redirect_) begin
        num$write_data = (head_tail_delta == 0) ? max_entries : { { 5-4 { 1'b0 } }, head_tail_delta };
      end
      else begin
        if ((register_success^commit_call)) begin
          if (register_success) begin
            num$write_data = (num$read_data+1);
          end
          else begin
            if (commit_call) begin
              num$write_data = (num$read_data-1);
            end
            else begin
            end
          end
        end
        else begin
        end
      end
    end
  end


endmodule // ControlFlowManager_0x734ebf4161405225

//-----------------------------------------------------------------------------
// Register_0x5d4baebedb8e9d8
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(4)); write <C> (data: Bits(4)) -> ()", "reset_value": 0}
// PyMTL: verilator_xinit = zeros
module Register_0x5d4baebedb8e9d8
(
  input  logic [   0:0] clk,
  output logic [   3:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [   3:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [   3:0] reg_value;

  // localparam declarations
  localparam reset_value = 0;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.reset:
  //           s.reg_value.n = reset_value
  //         elif s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      reg_value <= reset_value;
    end
    else begin
      if (update) begin
        reg_value <= write_data;
      end
      else begin
      end
    end
  end


endmodule // Register_0x5d4baebedb8e9d8

//-----------------------------------------------------------------------------
// OneHotEncoder_0x6ddac805079c9f17
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.onehot {"enable": true, "noutbits": 2}
// PyMTL: verilator_xinit = zeros
module OneHotEncoder_0x6ddac805079c9f17
(
  input  logic [   0:0] clk,
  input  logic [   0:0] encode_call,
  input  logic [   0:0] encode_number,
  output logic  [   1:0] encode_onehot,
  input  logic [   0:0] reset
);



  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[0] = (encode_call&&(encode_number == 0));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[1] = (encode_call&&(encode_number == 1));
  end


endmodule // OneHotEncoder_0x6ddac805079c9f17

//-----------------------------------------------------------------------------
// Register_0xae4a367f21f784a
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(5)); write <C> (data: Bits(5)) -> ()", "reset_value": 0}
// PyMTL: verilator_xinit = zeros
module Register_0xae4a367f21f784a
(
  input  logic [   0:0] clk,
  output logic [   4:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [   4:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [   4:0] reg_value;

  // localparam declarations
  localparam reset_value = 0;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.reset:
  //           s.reg_value.n = reset_value
  //         elif s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      reg_value <= reset_value;
    end
    else begin
      if (update) begin
        reg_value <= write_data;
      end
      else begin
      end
    end
  end


endmodule // Register_0xae4a367f21f784a

//-----------------------------------------------------------------------------
// AsynchronousRAM_0x7bb0942938a43a9
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.async_ram {"interface": "read[1] (addr: Bits(1)) -> (data: Bits(64)); write[1] <C> (data: Bits(64), addr: Bits(1)) -> ()", "reset_values": null}
// PyMTL: verilator_xinit = zeros
module AsynchronousRAM_0x7bb0942938a43a9
(
  input  logic [   0:0] clk,
  input  logic [   0:0] read_addr$000,
  output logic [  63:0] read_data$000,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_addr$000,
  input  logic [   0:0] write_call$000,
  input  logic [  63:0] write_data$000
);

  // logic declarations
  logic   [  63:0] regs$000;
  logic   [  63:0] regs$001;


  // localparam declarations
  localparam num_read_ports = 1;
  localparam num_write_ports = 1;

  // loop variable declarations
  integer i;


  // array declarations
  logic   [   0:0] read_addr[0:0];
  assign read_addr[  0] = read_addr$000;
  logic    [  63:0] read_data[0:0];
  assign read_data$000 = read_data[  0];
  logic    [  63:0] regs[0:1];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  logic   [   0:0] write_addr[0:0];
  assign write_addr[  0] = write_addr$000;
  logic   [   0:0] write_call[0:0];
  assign write_call[  0] = write_call$000;
  logic   [  63:0] write_data[0:0];
  assign write_data[  0] = write_data$000;

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def handle_writes():
  //         for i in range(num_write_ports):
  //           if s.write_call[i]:
  //             s.regs[s.write_addr[i]].n = s.write_data[i]

  // logic for handle_writes()
  always @ (posedge clk) begin
    for (i=0; i < num_write_ports; i=i+1)
    begin
      if (write_call[i]) begin
        regs[write_addr[i]] <= write_data[i];
      end
      else begin
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_reads():
  //         for i in range(num_read_ports):
  //           s.read_data[i].v = s.regs[s.read_addr[i]]

  // logic for handle_reads()
  always @ (*) begin
    for (i=0; i < num_read_ports; i=i+1)
    begin
      read_data[i] = regs[read_addr[i]];
    end
  end


endmodule // AsynchronousRAM_0x7bb0942938a43a9

//-----------------------------------------------------------------------------
// Register_0x19ffe7c045ca5b3a
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(1)); write <C> (data: Bits(1)) -> ()", "reset_value": 0}
// PyMTL: verilator_xinit = zeros
module Register_0x19ffe7c045ca5b3a
(
  input  logic [   0:0] clk,
  output logic [   0:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [   0:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [   0:0] reg_value;

  // localparam declarations
  localparam reset_value = 0;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.reset:
  //           s.reg_value.n = reset_value
  //         elif s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      reg_value <= reset_value;
    end
    else begin
      if (update) begin
        reg_value <= write_data;
      end
      else begin
      end
    end
  end


endmodule // Register_0x19ffe7c045ca5b3a

//-----------------------------------------------------------------------------
// Register_0x60b9ec19bb3fa768
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(2)); write <C> (data: Bits(2)) -> ()", "reset_value": 0}
// PyMTL: verilator_xinit = zeros
module Register_0x60b9ec19bb3fa768
(
  input  logic [   0:0] clk,
  output logic [   1:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [   1:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [   1:0] reg_value;

  // localparam declarations
  localparam reset_value = 0;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.reset:
  //           s.reg_value.n = reset_value
  //         elif s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      reg_value <= reset_value;
    end
    else begin
      if (update) begin
        reg_value <= write_data;
      end
      else begin
      end
    end
  end


endmodule // Register_0x60b9ec19bb3fa768

//-----------------------------------------------------------------------------
// Commit_0x7d8cae7cdd7a2d86
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.backend.commit {"interface": "kill_notify (msg: Bits(5)) -> ()", "rob_size": 16}
// PyMTL: verilator_xinit = zeros
module Commit_0x7d8cae7cdd7a2d86
(
  output logic [   0:0] cflow_commit_call,
  output logic [   1:0] cflow_commit_status,
  input  logic [   0:0] cflow_get_head_rdy,
  input  logic [   3:0] cflow_get_head_seq,
  input  logic [   0:0] clk,
  output logic  [   0:0] dataflow_commit_call,
  output logic  [   5:0] dataflow_commit_tag,
  input  logic [ 141:0] in_peek_msg,
  input  logic [   0:0] in_peek_rdy,
  output logic [   0:0] in_take_call,
  input  logic [   4:0] kill_notify_msg,
  input  logic [   0:0] reset
);

  // logic declarations
  logic   [   0:0] advance;
  logic   [   3:0] seq_num;


  // register declarations
  logic    [   0:0] rob_remove;

  // localparam declarations
  localparam PIPELINE_MSG_STATUS_VALID = 2'd0;

  // rob temporaries
  logic   [   3:0] rob$check_done_idx;
  logic   [   0:0] rob$clk;
  logic   [   0:0] rob$free_call;
  logic   [   4:0] rob$kill_notify_msg;
  logic   [   3:0] rob$free_idx;
  logic   [ 141:0] rob$add_value;
  logic   [   0:0] rob$reset;
  logic   [   0:0] rob$add_call;
  logic   [   3:0] rob$add_idx;
  logic   [   1:0] rob$add_kill_opaque;
  logic   [ 141:0] rob$free_value;
  logic   [   0:0] rob$check_done_is_rdy;

  ReorderBuffer_0x46a5141874a5c0a2 rob
  (
    .check_done_idx    ( rob$check_done_idx ),
    .clk               ( rob$clk ),
    .free_call         ( rob$free_call ),
    .kill_notify_msg   ( rob$kill_notify_msg ),
    .free_idx          ( rob$free_idx ),
    .add_value         ( rob$add_value ),
    .reset             ( rob$reset ),
    .add_call          ( rob$add_call ),
    .add_idx           ( rob$add_idx ),
    .add_kill_opaque   ( rob$add_kill_opaque ),
    .free_value        ( rob$free_value ),
    .check_done_is_rdy ( rob$check_done_is_rdy )
  );

  // signal connections
  assign advance             = in_peek_rdy;
  assign cflow_commit_call   = rob_remove;
  assign cflow_commit_status = rob$free_value[1:0];
  assign in_take_call        = advance;
  assign rob$add_call        = advance;
  assign rob$add_idx         = seq_num;
  assign rob$add_value       = in_peek_msg;
  assign rob$check_done_idx  = cflow_get_head_seq;
  assign rob$clk             = clk;
  assign rob$free_call       = rob_remove;
  assign rob$free_idx        = cflow_get_head_seq;
  assign rob$kill_notify_msg = kill_notify_msg;
  assign rob$reset           = reset;
  assign seq_num             = in_peek_msg[69:66];


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def set_rob_remove():
  //       s.rob_remove.v = s.cflow_get_head_rdy and s.rob.check_done_is_rdy

  // logic for set_rob_remove()
  always @ (*) begin
    rob_remove = (cflow_get_head_rdy&&rob$check_done_is_rdy);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_commit():
  //       s.dataflow_commit_call.v = 0
  //       s.dataflow_commit_tag.v = 0
  //
  //       # The head is ready to commit
  //       if s.rob_remove:
  //         if s.rob.free_value.hdr_status == PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID:
  //           if s.rob.free_value.rd_val:
  //             s.dataflow_commit_call.v = 1
  //             s.dataflow_commit_tag.v = s.rob.free_value.rd
  //         else:
  //           # TODO handle exception
  //           # PYMTL_BROKEN pass doesn't work
  //           # pass
  //           s.dataflow_commit_tag.v = 0

  // logic for handle_commit()
  always @ (*) begin
    dataflow_commit_call = 0;
    dataflow_commit_tag = 0;
    if (rob_remove) begin
      if ((rob$free_value[(2)-1:0] == PIPELINE_MSG_STATUS_VALID)) begin
        if (rob$free_value[(75)-1:74]) begin
          dataflow_commit_call = 1;
          dataflow_commit_tag = rob$free_value[(81)-1:75];
        end
        else begin
        end
      end
      else begin
        dataflow_commit_tag = 0;
      end
    end
    else begin
    end
  end


endmodule // Commit_0x7d8cae7cdd7a2d86

//-----------------------------------------------------------------------------
// ReorderBuffer_0x46a5141874a5c0a2
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.reorder_buffer {"interface": "add <C> (kill_opaque: Bits(2), idx: Bits(4), value: Bits(142)) -> (); check_done (idx: Bits(4)) -> (is_rdy: Bits(1)); free <C> (idx: Bits(4)) -> (value: Bits(142)); kill_notify (msg: Bits(5)) -> ()", "make_kill": "<function make_kill at 0x7f0068be79b0>"}
// PyMTL: verilator_xinit = zeros
module ReorderBuffer_0x46a5141874a5c0a2
(
  input  logic [   0:0] add_call,
  input  logic [   3:0] add_idx,
  input  logic [   1:0] add_kill_opaque,
  input  logic [ 141:0] add_value,
  input  logic [   3:0] check_done_idx,
  output logic [   0:0] check_done_is_rdy,
  input  logic [   0:0] clk,
  input  logic [   0:0] free_call,
  input  logic [   3:0] free_idx,
  output logic [ 141:0] free_value,
  input  logic [   4:0] kill_notify_msg,
  input  logic [   0:0] reset
);

  // valids_$000 temporaries
  logic   [   4:0] valids_$000$kill_notify_msg;
  logic   [   0:0] valids_$000$clk;
  logic   [   1:0] valids_$000$add_msg;
  logic   [   0:0] valids_$000$reset;
  logic   [   0:0] valids_$000$add_call;
  logic   [   0:0] valids_$000$take_call;
  logic   [   1:0] valids_$000$peek_msg;
  logic   [   0:0] valids_$000$add_rdy;
  logic   [   0:0] valids_$000$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$000
  (
    .kill_notify_msg ( valids_$000$kill_notify_msg ),
    .clk             ( valids_$000$clk ),
    .add_msg         ( valids_$000$add_msg ),
    .reset           ( valids_$000$reset ),
    .add_call        ( valids_$000$add_call ),
    .take_call       ( valids_$000$take_call ),
    .peek_msg        ( valids_$000$peek_msg ),
    .add_rdy         ( valids_$000$add_rdy ),
    .peek_rdy        ( valids_$000$peek_rdy )
  );

  // valids_$001 temporaries
  logic   [   4:0] valids_$001$kill_notify_msg;
  logic   [   0:0] valids_$001$clk;
  logic   [   1:0] valids_$001$add_msg;
  logic   [   0:0] valids_$001$reset;
  logic   [   0:0] valids_$001$add_call;
  logic   [   0:0] valids_$001$take_call;
  logic   [   1:0] valids_$001$peek_msg;
  logic   [   0:0] valids_$001$add_rdy;
  logic   [   0:0] valids_$001$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$001
  (
    .kill_notify_msg ( valids_$001$kill_notify_msg ),
    .clk             ( valids_$001$clk ),
    .add_msg         ( valids_$001$add_msg ),
    .reset           ( valids_$001$reset ),
    .add_call        ( valids_$001$add_call ),
    .take_call       ( valids_$001$take_call ),
    .peek_msg        ( valids_$001$peek_msg ),
    .add_rdy         ( valids_$001$add_rdy ),
    .peek_rdy        ( valids_$001$peek_rdy )
  );

  // valids_$002 temporaries
  logic   [   4:0] valids_$002$kill_notify_msg;
  logic   [   0:0] valids_$002$clk;
  logic   [   1:0] valids_$002$add_msg;
  logic   [   0:0] valids_$002$reset;
  logic   [   0:0] valids_$002$add_call;
  logic   [   0:0] valids_$002$take_call;
  logic   [   1:0] valids_$002$peek_msg;
  logic   [   0:0] valids_$002$add_rdy;
  logic   [   0:0] valids_$002$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$002
  (
    .kill_notify_msg ( valids_$002$kill_notify_msg ),
    .clk             ( valids_$002$clk ),
    .add_msg         ( valids_$002$add_msg ),
    .reset           ( valids_$002$reset ),
    .add_call        ( valids_$002$add_call ),
    .take_call       ( valids_$002$take_call ),
    .peek_msg        ( valids_$002$peek_msg ),
    .add_rdy         ( valids_$002$add_rdy ),
    .peek_rdy        ( valids_$002$peek_rdy )
  );

  // valids_$003 temporaries
  logic   [   4:0] valids_$003$kill_notify_msg;
  logic   [   0:0] valids_$003$clk;
  logic   [   1:0] valids_$003$add_msg;
  logic   [   0:0] valids_$003$reset;
  logic   [   0:0] valids_$003$add_call;
  logic   [   0:0] valids_$003$take_call;
  logic   [   1:0] valids_$003$peek_msg;
  logic   [   0:0] valids_$003$add_rdy;
  logic   [   0:0] valids_$003$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$003
  (
    .kill_notify_msg ( valids_$003$kill_notify_msg ),
    .clk             ( valids_$003$clk ),
    .add_msg         ( valids_$003$add_msg ),
    .reset           ( valids_$003$reset ),
    .add_call        ( valids_$003$add_call ),
    .take_call       ( valids_$003$take_call ),
    .peek_msg        ( valids_$003$peek_msg ),
    .add_rdy         ( valids_$003$add_rdy ),
    .peek_rdy        ( valids_$003$peek_rdy )
  );

  // valids_$004 temporaries
  logic   [   4:0] valids_$004$kill_notify_msg;
  logic   [   0:0] valids_$004$clk;
  logic   [   1:0] valids_$004$add_msg;
  logic   [   0:0] valids_$004$reset;
  logic   [   0:0] valids_$004$add_call;
  logic   [   0:0] valids_$004$take_call;
  logic   [   1:0] valids_$004$peek_msg;
  logic   [   0:0] valids_$004$add_rdy;
  logic   [   0:0] valids_$004$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$004
  (
    .kill_notify_msg ( valids_$004$kill_notify_msg ),
    .clk             ( valids_$004$clk ),
    .add_msg         ( valids_$004$add_msg ),
    .reset           ( valids_$004$reset ),
    .add_call        ( valids_$004$add_call ),
    .take_call       ( valids_$004$take_call ),
    .peek_msg        ( valids_$004$peek_msg ),
    .add_rdy         ( valids_$004$add_rdy ),
    .peek_rdy        ( valids_$004$peek_rdy )
  );

  // valids_$005 temporaries
  logic   [   4:0] valids_$005$kill_notify_msg;
  logic   [   0:0] valids_$005$clk;
  logic   [   1:0] valids_$005$add_msg;
  logic   [   0:0] valids_$005$reset;
  logic   [   0:0] valids_$005$add_call;
  logic   [   0:0] valids_$005$take_call;
  logic   [   1:0] valids_$005$peek_msg;
  logic   [   0:0] valids_$005$add_rdy;
  logic   [   0:0] valids_$005$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$005
  (
    .kill_notify_msg ( valids_$005$kill_notify_msg ),
    .clk             ( valids_$005$clk ),
    .add_msg         ( valids_$005$add_msg ),
    .reset           ( valids_$005$reset ),
    .add_call        ( valids_$005$add_call ),
    .take_call       ( valids_$005$take_call ),
    .peek_msg        ( valids_$005$peek_msg ),
    .add_rdy         ( valids_$005$add_rdy ),
    .peek_rdy        ( valids_$005$peek_rdy )
  );

  // valids_$006 temporaries
  logic   [   4:0] valids_$006$kill_notify_msg;
  logic   [   0:0] valids_$006$clk;
  logic   [   1:0] valids_$006$add_msg;
  logic   [   0:0] valids_$006$reset;
  logic   [   0:0] valids_$006$add_call;
  logic   [   0:0] valids_$006$take_call;
  logic   [   1:0] valids_$006$peek_msg;
  logic   [   0:0] valids_$006$add_rdy;
  logic   [   0:0] valids_$006$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$006
  (
    .kill_notify_msg ( valids_$006$kill_notify_msg ),
    .clk             ( valids_$006$clk ),
    .add_msg         ( valids_$006$add_msg ),
    .reset           ( valids_$006$reset ),
    .add_call        ( valids_$006$add_call ),
    .take_call       ( valids_$006$take_call ),
    .peek_msg        ( valids_$006$peek_msg ),
    .add_rdy         ( valids_$006$add_rdy ),
    .peek_rdy        ( valids_$006$peek_rdy )
  );

  // valids_$007 temporaries
  logic   [   4:0] valids_$007$kill_notify_msg;
  logic   [   0:0] valids_$007$clk;
  logic   [   1:0] valids_$007$add_msg;
  logic   [   0:0] valids_$007$reset;
  logic   [   0:0] valids_$007$add_call;
  logic   [   0:0] valids_$007$take_call;
  logic   [   1:0] valids_$007$peek_msg;
  logic   [   0:0] valids_$007$add_rdy;
  logic   [   0:0] valids_$007$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$007
  (
    .kill_notify_msg ( valids_$007$kill_notify_msg ),
    .clk             ( valids_$007$clk ),
    .add_msg         ( valids_$007$add_msg ),
    .reset           ( valids_$007$reset ),
    .add_call        ( valids_$007$add_call ),
    .take_call       ( valids_$007$take_call ),
    .peek_msg        ( valids_$007$peek_msg ),
    .add_rdy         ( valids_$007$add_rdy ),
    .peek_rdy        ( valids_$007$peek_rdy )
  );

  // valids_$008 temporaries
  logic   [   4:0] valids_$008$kill_notify_msg;
  logic   [   0:0] valids_$008$clk;
  logic   [   1:0] valids_$008$add_msg;
  logic   [   0:0] valids_$008$reset;
  logic   [   0:0] valids_$008$add_call;
  logic   [   0:0] valids_$008$take_call;
  logic   [   1:0] valids_$008$peek_msg;
  logic   [   0:0] valids_$008$add_rdy;
  logic   [   0:0] valids_$008$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$008
  (
    .kill_notify_msg ( valids_$008$kill_notify_msg ),
    .clk             ( valids_$008$clk ),
    .add_msg         ( valids_$008$add_msg ),
    .reset           ( valids_$008$reset ),
    .add_call        ( valids_$008$add_call ),
    .take_call       ( valids_$008$take_call ),
    .peek_msg        ( valids_$008$peek_msg ),
    .add_rdy         ( valids_$008$add_rdy ),
    .peek_rdy        ( valids_$008$peek_rdy )
  );

  // valids_$009 temporaries
  logic   [   4:0] valids_$009$kill_notify_msg;
  logic   [   0:0] valids_$009$clk;
  logic   [   1:0] valids_$009$add_msg;
  logic   [   0:0] valids_$009$reset;
  logic   [   0:0] valids_$009$add_call;
  logic   [   0:0] valids_$009$take_call;
  logic   [   1:0] valids_$009$peek_msg;
  logic   [   0:0] valids_$009$add_rdy;
  logic   [   0:0] valids_$009$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$009
  (
    .kill_notify_msg ( valids_$009$kill_notify_msg ),
    .clk             ( valids_$009$clk ),
    .add_msg         ( valids_$009$add_msg ),
    .reset           ( valids_$009$reset ),
    .add_call        ( valids_$009$add_call ),
    .take_call       ( valids_$009$take_call ),
    .peek_msg        ( valids_$009$peek_msg ),
    .add_rdy         ( valids_$009$add_rdy ),
    .peek_rdy        ( valids_$009$peek_rdy )
  );

  // valids_$010 temporaries
  logic   [   4:0] valids_$010$kill_notify_msg;
  logic   [   0:0] valids_$010$clk;
  logic   [   1:0] valids_$010$add_msg;
  logic   [   0:0] valids_$010$reset;
  logic   [   0:0] valids_$010$add_call;
  logic   [   0:0] valids_$010$take_call;
  logic   [   1:0] valids_$010$peek_msg;
  logic   [   0:0] valids_$010$add_rdy;
  logic   [   0:0] valids_$010$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$010
  (
    .kill_notify_msg ( valids_$010$kill_notify_msg ),
    .clk             ( valids_$010$clk ),
    .add_msg         ( valids_$010$add_msg ),
    .reset           ( valids_$010$reset ),
    .add_call        ( valids_$010$add_call ),
    .take_call       ( valids_$010$take_call ),
    .peek_msg        ( valids_$010$peek_msg ),
    .add_rdy         ( valids_$010$add_rdy ),
    .peek_rdy        ( valids_$010$peek_rdy )
  );

  // valids_$011 temporaries
  logic   [   4:0] valids_$011$kill_notify_msg;
  logic   [   0:0] valids_$011$clk;
  logic   [   1:0] valids_$011$add_msg;
  logic   [   0:0] valids_$011$reset;
  logic   [   0:0] valids_$011$add_call;
  logic   [   0:0] valids_$011$take_call;
  logic   [   1:0] valids_$011$peek_msg;
  logic   [   0:0] valids_$011$add_rdy;
  logic   [   0:0] valids_$011$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$011
  (
    .kill_notify_msg ( valids_$011$kill_notify_msg ),
    .clk             ( valids_$011$clk ),
    .add_msg         ( valids_$011$add_msg ),
    .reset           ( valids_$011$reset ),
    .add_call        ( valids_$011$add_call ),
    .take_call       ( valids_$011$take_call ),
    .peek_msg        ( valids_$011$peek_msg ),
    .add_rdy         ( valids_$011$add_rdy ),
    .peek_rdy        ( valids_$011$peek_rdy )
  );

  // valids_$012 temporaries
  logic   [   4:0] valids_$012$kill_notify_msg;
  logic   [   0:0] valids_$012$clk;
  logic   [   1:0] valids_$012$add_msg;
  logic   [   0:0] valids_$012$reset;
  logic   [   0:0] valids_$012$add_call;
  logic   [   0:0] valids_$012$take_call;
  logic   [   1:0] valids_$012$peek_msg;
  logic   [   0:0] valids_$012$add_rdy;
  logic   [   0:0] valids_$012$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$012
  (
    .kill_notify_msg ( valids_$012$kill_notify_msg ),
    .clk             ( valids_$012$clk ),
    .add_msg         ( valids_$012$add_msg ),
    .reset           ( valids_$012$reset ),
    .add_call        ( valids_$012$add_call ),
    .take_call       ( valids_$012$take_call ),
    .peek_msg        ( valids_$012$peek_msg ),
    .add_rdy         ( valids_$012$add_rdy ),
    .peek_rdy        ( valids_$012$peek_rdy )
  );

  // valids_$013 temporaries
  logic   [   4:0] valids_$013$kill_notify_msg;
  logic   [   0:0] valids_$013$clk;
  logic   [   1:0] valids_$013$add_msg;
  logic   [   0:0] valids_$013$reset;
  logic   [   0:0] valids_$013$add_call;
  logic   [   0:0] valids_$013$take_call;
  logic   [   1:0] valids_$013$peek_msg;
  logic   [   0:0] valids_$013$add_rdy;
  logic   [   0:0] valids_$013$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$013
  (
    .kill_notify_msg ( valids_$013$kill_notify_msg ),
    .clk             ( valids_$013$clk ),
    .add_msg         ( valids_$013$add_msg ),
    .reset           ( valids_$013$reset ),
    .add_call        ( valids_$013$add_call ),
    .take_call       ( valids_$013$take_call ),
    .peek_msg        ( valids_$013$peek_msg ),
    .add_rdy         ( valids_$013$add_rdy ),
    .peek_rdy        ( valids_$013$peek_rdy )
  );

  // valids_$014 temporaries
  logic   [   4:0] valids_$014$kill_notify_msg;
  logic   [   0:0] valids_$014$clk;
  logic   [   1:0] valids_$014$add_msg;
  logic   [   0:0] valids_$014$reset;
  logic   [   0:0] valids_$014$add_call;
  logic   [   0:0] valids_$014$take_call;
  logic   [   1:0] valids_$014$peek_msg;
  logic   [   0:0] valids_$014$add_rdy;
  logic   [   0:0] valids_$014$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$014
  (
    .kill_notify_msg ( valids_$014$kill_notify_msg ),
    .clk             ( valids_$014$clk ),
    .add_msg         ( valids_$014$add_msg ),
    .reset           ( valids_$014$reset ),
    .add_call        ( valids_$014$add_call ),
    .take_call       ( valids_$014$take_call ),
    .peek_msg        ( valids_$014$peek_msg ),
    .add_rdy         ( valids_$014$add_rdy ),
    .peek_rdy        ( valids_$014$peek_rdy )
  );

  // valids_$015 temporaries
  logic   [   4:0] valids_$015$kill_notify_msg;
  logic   [   0:0] valids_$015$clk;
  logic   [   1:0] valids_$015$add_msg;
  logic   [   0:0] valids_$015$reset;
  logic   [   0:0] valids_$015$add_call;
  logic   [   0:0] valids_$015$take_call;
  logic   [   1:0] valids_$015$peek_msg;
  logic   [   0:0] valids_$015$add_rdy;
  logic   [   0:0] valids_$015$peek_rdy;

  GenValidValueManager9Lmake_kill_0x70f4a78affa17bfb valids_$015
  (
    .kill_notify_msg ( valids_$015$kill_notify_msg ),
    .clk             ( valids_$015$clk ),
    .add_msg         ( valids_$015$add_msg ),
    .reset           ( valids_$015$reset ),
    .add_call        ( valids_$015$add_call ),
    .take_call       ( valids_$015$take_call ),
    .peek_msg        ( valids_$015$peek_msg ),
    .add_rdy         ( valids_$015$add_rdy ),
    .peek_rdy        ( valids_$015$peek_rdy )
  );

  // add_encoder_ temporaries
  logic   [   0:0] add_encoder_$encode_call;
  logic   [   0:0] add_encoder_$clk;
  logic   [   0:0] add_encoder_$reset;
  logic   [   3:0] add_encoder_$encode_number;
  logic   [  15:0] add_encoder_$encode_onehot;

  OneHotEncoder_0x1fe0e9741db02a15 add_encoder_
  (
    .encode_call   ( add_encoder_$encode_call ),
    .clk           ( add_encoder_$clk ),
    .reset         ( add_encoder_$reset ),
    .encode_number ( add_encoder_$encode_number ),
    .encode_onehot ( add_encoder_$encode_onehot )
  );

  // free_encoder_ temporaries
  logic   [   0:0] free_encoder_$encode_call;
  logic   [   0:0] free_encoder_$clk;
  logic   [   0:0] free_encoder_$reset;
  logic   [   3:0] free_encoder_$encode_number;
  logic   [  15:0] free_encoder_$encode_onehot;

  OneHotEncoder_0x1fe0e9741db02a15 free_encoder_
  (
    .encode_call   ( free_encoder_$encode_call ),
    .clk           ( free_encoder_$clk ),
    .reset         ( free_encoder_$reset ),
    .encode_number ( free_encoder_$encode_number ),
    .encode_onehot ( free_encoder_$encode_onehot )
  );

  // entries_ temporaries
  logic   [   0:0] entries_$clk;
  logic   [   3:0] entries_$write_addr$000;
  logic   [   3:0] entries_$read_addr$000;
  logic   [   0:0] entries_$write_call$000;
  logic   [ 141:0] entries_$write_data$000;
  logic   [   0:0] entries_$reset;
  logic   [ 141:0] entries_$read_data$000;

  AsynchronousRAM_0x3c5ad87dd535d6cd entries_
  (
    .clk            ( entries_$clk ),
    .write_addr$000 ( entries_$write_addr$000 ),
    .read_addr$000  ( entries_$read_addr$000 ),
    .write_call$000 ( entries_$write_call$000 ),
    .write_data$000 ( entries_$write_data$000 ),
    .reset          ( entries_$reset ),
    .read_data$000  ( entries_$read_data$000 )
  );

  // mux_done_ temporaries
  logic   [   0:0] mux_done_$mux_in_$000;
  logic   [   0:0] mux_done_$mux_in_$001;
  logic   [   0:0] mux_done_$mux_in_$002;
  logic   [   0:0] mux_done_$mux_in_$003;
  logic   [   0:0] mux_done_$mux_in_$004;
  logic   [   0:0] mux_done_$mux_in_$005;
  logic   [   0:0] mux_done_$mux_in_$006;
  logic   [   0:0] mux_done_$mux_in_$007;
  logic   [   0:0] mux_done_$mux_in_$008;
  logic   [   0:0] mux_done_$mux_in_$009;
  logic   [   0:0] mux_done_$mux_in_$010;
  logic   [   0:0] mux_done_$mux_in_$011;
  logic   [   0:0] mux_done_$mux_in_$012;
  logic   [   0:0] mux_done_$mux_in_$013;
  logic   [   0:0] mux_done_$mux_in_$014;
  logic   [   0:0] mux_done_$mux_in_$015;
  logic   [   0:0] mux_done_$clk;
  logic   [   0:0] mux_done_$reset;
  logic   [   3:0] mux_done_$mux_select;
  logic   [   0:0] mux_done_$mux_out;

  Mux_0x71ecd1c0a6217ee5 mux_done_
  (
    .mux_in_$000 ( mux_done_$mux_in_$000 ),
    .mux_in_$001 ( mux_done_$mux_in_$001 ),
    .mux_in_$002 ( mux_done_$mux_in_$002 ),
    .mux_in_$003 ( mux_done_$mux_in_$003 ),
    .mux_in_$004 ( mux_done_$mux_in_$004 ),
    .mux_in_$005 ( mux_done_$mux_in_$005 ),
    .mux_in_$006 ( mux_done_$mux_in_$006 ),
    .mux_in_$007 ( mux_done_$mux_in_$007 ),
    .mux_in_$008 ( mux_done_$mux_in_$008 ),
    .mux_in_$009 ( mux_done_$mux_in_$009 ),
    .mux_in_$010 ( mux_done_$mux_in_$010 ),
    .mux_in_$011 ( mux_done_$mux_in_$011 ),
    .mux_in_$012 ( mux_done_$mux_in_$012 ),
    .mux_in_$013 ( mux_done_$mux_in_$013 ),
    .mux_in_$014 ( mux_done_$mux_in_$014 ),
    .mux_in_$015 ( mux_done_$mux_in_$015 ),
    .clk         ( mux_done_$clk ),
    .reset       ( mux_done_$reset ),
    .mux_select  ( mux_done_$mux_select ),
    .mux_out     ( mux_done_$mux_out )
  );

  // signal connections
  assign add_encoder_$clk            = clk;
  assign add_encoder_$encode_call    = add_call;
  assign add_encoder_$encode_number  = add_idx;
  assign add_encoder_$reset          = reset;
  assign check_done_is_rdy           = mux_done_$mux_out;
  assign entries_$clk                = clk;
  assign entries_$read_addr$000      = free_idx;
  assign entries_$reset              = reset;
  assign entries_$write_addr$000     = add_idx;
  assign entries_$write_call$000     = add_call;
  assign entries_$write_data$000     = add_value;
  assign free_encoder_$clk           = clk;
  assign free_encoder_$encode_call   = free_call;
  assign free_encoder_$encode_number = free_idx;
  assign free_encoder_$reset         = reset;
  assign free_value                  = entries_$read_data$000;
  assign mux_done_$clk               = clk;
  assign mux_done_$mux_in_$000       = valids_$000$peek_rdy;
  assign mux_done_$mux_in_$001       = valids_$001$peek_rdy;
  assign mux_done_$mux_in_$002       = valids_$002$peek_rdy;
  assign mux_done_$mux_in_$003       = valids_$003$peek_rdy;
  assign mux_done_$mux_in_$004       = valids_$004$peek_rdy;
  assign mux_done_$mux_in_$005       = valids_$005$peek_rdy;
  assign mux_done_$mux_in_$006       = valids_$006$peek_rdy;
  assign mux_done_$mux_in_$007       = valids_$007$peek_rdy;
  assign mux_done_$mux_in_$008       = valids_$008$peek_rdy;
  assign mux_done_$mux_in_$009       = valids_$009$peek_rdy;
  assign mux_done_$mux_in_$010       = valids_$010$peek_rdy;
  assign mux_done_$mux_in_$011       = valids_$011$peek_rdy;
  assign mux_done_$mux_in_$012       = valids_$012$peek_rdy;
  assign mux_done_$mux_in_$013       = valids_$013$peek_rdy;
  assign mux_done_$mux_in_$014       = valids_$014$peek_rdy;
  assign mux_done_$mux_in_$015       = valids_$015$peek_rdy;
  assign mux_done_$mux_select        = check_done_idx;
  assign mux_done_$reset             = reset;
  assign valids_$000$add_call        = add_encoder_$encode_onehot[0];
  assign valids_$000$add_msg         = add_kill_opaque;
  assign valids_$000$clk             = clk;
  assign valids_$000$kill_notify_msg = kill_notify_msg;
  assign valids_$000$reset           = reset;
  assign valids_$000$take_call       = free_encoder_$encode_onehot[0];
  assign valids_$001$add_call        = add_encoder_$encode_onehot[1];
  assign valids_$001$add_msg         = add_kill_opaque;
  assign valids_$001$clk             = clk;
  assign valids_$001$kill_notify_msg = kill_notify_msg;
  assign valids_$001$reset           = reset;
  assign valids_$001$take_call       = free_encoder_$encode_onehot[1];
  assign valids_$002$add_call        = add_encoder_$encode_onehot[2];
  assign valids_$002$add_msg         = add_kill_opaque;
  assign valids_$002$clk             = clk;
  assign valids_$002$kill_notify_msg = kill_notify_msg;
  assign valids_$002$reset           = reset;
  assign valids_$002$take_call       = free_encoder_$encode_onehot[2];
  assign valids_$003$add_call        = add_encoder_$encode_onehot[3];
  assign valids_$003$add_msg         = add_kill_opaque;
  assign valids_$003$clk             = clk;
  assign valids_$003$kill_notify_msg = kill_notify_msg;
  assign valids_$003$reset           = reset;
  assign valids_$003$take_call       = free_encoder_$encode_onehot[3];
  assign valids_$004$add_call        = add_encoder_$encode_onehot[4];
  assign valids_$004$add_msg         = add_kill_opaque;
  assign valids_$004$clk             = clk;
  assign valids_$004$kill_notify_msg = kill_notify_msg;
  assign valids_$004$reset           = reset;
  assign valids_$004$take_call       = free_encoder_$encode_onehot[4];
  assign valids_$005$add_call        = add_encoder_$encode_onehot[5];
  assign valids_$005$add_msg         = add_kill_opaque;
  assign valids_$005$clk             = clk;
  assign valids_$005$kill_notify_msg = kill_notify_msg;
  assign valids_$005$reset           = reset;
  assign valids_$005$take_call       = free_encoder_$encode_onehot[5];
  assign valids_$006$add_call        = add_encoder_$encode_onehot[6];
  assign valids_$006$add_msg         = add_kill_opaque;
  assign valids_$006$clk             = clk;
  assign valids_$006$kill_notify_msg = kill_notify_msg;
  assign valids_$006$reset           = reset;
  assign valids_$006$take_call       = free_encoder_$encode_onehot[6];
  assign valids_$007$add_call        = add_encoder_$encode_onehot[7];
  assign valids_$007$add_msg         = add_kill_opaque;
  assign valids_$007$clk             = clk;
  assign valids_$007$kill_notify_msg = kill_notify_msg;
  assign valids_$007$reset           = reset;
  assign valids_$007$take_call       = free_encoder_$encode_onehot[7];
  assign valids_$008$add_call        = add_encoder_$encode_onehot[8];
  assign valids_$008$add_msg         = add_kill_opaque;
  assign valids_$008$clk             = clk;
  assign valids_$008$kill_notify_msg = kill_notify_msg;
  assign valids_$008$reset           = reset;
  assign valids_$008$take_call       = free_encoder_$encode_onehot[8];
  assign valids_$009$add_call        = add_encoder_$encode_onehot[9];
  assign valids_$009$add_msg         = add_kill_opaque;
  assign valids_$009$clk             = clk;
  assign valids_$009$kill_notify_msg = kill_notify_msg;
  assign valids_$009$reset           = reset;
  assign valids_$009$take_call       = free_encoder_$encode_onehot[9];
  assign valids_$010$add_call        = add_encoder_$encode_onehot[10];
  assign valids_$010$add_msg         = add_kill_opaque;
  assign valids_$010$clk             = clk;
  assign valids_$010$kill_notify_msg = kill_notify_msg;
  assign valids_$010$reset           = reset;
  assign valids_$010$take_call       = free_encoder_$encode_onehot[10];
  assign valids_$011$add_call        = add_encoder_$encode_onehot[11];
  assign valids_$011$add_msg         = add_kill_opaque;
  assign valids_$011$clk             = clk;
  assign valids_$011$kill_notify_msg = kill_notify_msg;
  assign valids_$011$reset           = reset;
  assign valids_$011$take_call       = free_encoder_$encode_onehot[11];
  assign valids_$012$add_call        = add_encoder_$encode_onehot[12];
  assign valids_$012$add_msg         = add_kill_opaque;
  assign valids_$012$clk             = clk;
  assign valids_$012$kill_notify_msg = kill_notify_msg;
  assign valids_$012$reset           = reset;
  assign valids_$012$take_call       = free_encoder_$encode_onehot[12];
  assign valids_$013$add_call        = add_encoder_$encode_onehot[13];
  assign valids_$013$add_msg         = add_kill_opaque;
  assign valids_$013$clk             = clk;
  assign valids_$013$kill_notify_msg = kill_notify_msg;
  assign valids_$013$reset           = reset;
  assign valids_$013$take_call       = free_encoder_$encode_onehot[13];
  assign valids_$014$add_call        = add_encoder_$encode_onehot[14];
  assign valids_$014$add_msg         = add_kill_opaque;
  assign valids_$014$clk             = clk;
  assign valids_$014$kill_notify_msg = kill_notify_msg;
  assign valids_$014$reset           = reset;
  assign valids_$014$take_call       = free_encoder_$encode_onehot[14];
  assign valids_$015$add_call        = add_encoder_$encode_onehot[15];
  assign valids_$015$add_msg         = add_kill_opaque;
  assign valids_$015$clk             = clk;
  assign valids_$015$kill_notify_msg = kill_notify_msg;
  assign valids_$015$reset           = reset;
  assign valids_$015$take_call       = free_encoder_$encode_onehot[15];



endmodule // ReorderBuffer_0x46a5141874a5c0a2

//-----------------------------------------------------------------------------
// OneHotEncoder_0x1fe0e9741db02a15
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.onehot {"enable": true, "noutbits": 16}
// PyMTL: verilator_xinit = zeros
module OneHotEncoder_0x1fe0e9741db02a15
(
  input  logic [   0:0] clk,
  input  logic [   0:0] encode_call,
  input  logic [   3:0] encode_number,
  output logic  [  15:0] encode_onehot,
  input  logic [   0:0] reset
);



  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[0] = (encode_call&&(encode_number == 0));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[1] = (encode_call&&(encode_number == 1));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[2] = (encode_call&&(encode_number == 2));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[3] = (encode_call&&(encode_number == 3));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[4] = (encode_call&&(encode_number == 4));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[5] = (encode_call&&(encode_number == 5));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[6] = (encode_call&&(encode_number == 6));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[7] = (encode_call&&(encode_number == 7));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[8] = (encode_call&&(encode_number == 8));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[9] = (encode_call&&(encode_number == 9));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[10] = (encode_call&&(encode_number == 10));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[11] = (encode_call&&(encode_number == 11));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[12] = (encode_call&&(encode_number == 12));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[13] = (encode_call&&(encode_number == 13));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[14] = (encode_call&&(encode_number == 14));
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_encode(i=i):
  //           s.encode_onehot[i].v = s.encode_call and (s.encode_number == i)

  // logic for handle_encode()
  always @ (*) begin
    encode_onehot[15] = (encode_call&&(encode_number == 15));
  end


endmodule // OneHotEncoder_0x1fe0e9741db02a15

//-----------------------------------------------------------------------------
// AsynchronousRAM_0x3c5ad87dd535d6cd
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.async_ram {"interface": "read[1] (addr: Bits(4)) -> (data: Bits(142)); write[1] <C> (data: Bits(142), addr: Bits(4)) -> ()", "reset_values": null}
// PyMTL: verilator_xinit = zeros
module AsynchronousRAM_0x3c5ad87dd535d6cd
(
  input  logic [   0:0] clk,
  input  logic [   3:0] read_addr$000,
  output logic [ 141:0] read_data$000,
  input  logic [   0:0] reset,
  input  logic [   3:0] write_addr$000,
  input  logic [   0:0] write_call$000,
  input  logic [ 141:0] write_data$000
);

  // logic declarations
  logic   [ 141:0] regs$000;
  logic   [ 141:0] regs$001;
  logic   [ 141:0] regs$002;
  logic   [ 141:0] regs$003;
  logic   [ 141:0] regs$004;
  logic   [ 141:0] regs$005;
  logic   [ 141:0] regs$006;
  logic   [ 141:0] regs$007;
  logic   [ 141:0] regs$008;
  logic   [ 141:0] regs$009;
  logic   [ 141:0] regs$010;
  logic   [ 141:0] regs$011;
  logic   [ 141:0] regs$012;
  logic   [ 141:0] regs$013;
  logic   [ 141:0] regs$014;
  logic   [ 141:0] regs$015;


  // localparam declarations
  localparam num_read_ports = 1;
  localparam num_write_ports = 1;

  // loop variable declarations
  integer i;


  // array declarations
  logic   [   3:0] read_addr[0:0];
  assign read_addr[  0] = read_addr$000;
  logic    [ 141:0] read_data[0:0];
  assign read_data$000 = read_data[  0];
  logic    [ 141:0] regs[0:15];
  assign regs$000 = regs[  0];
  assign regs$001 = regs[  1];
  assign regs$002 = regs[  2];
  assign regs$003 = regs[  3];
  assign regs$004 = regs[  4];
  assign regs$005 = regs[  5];
  assign regs$006 = regs[  6];
  assign regs$007 = regs[  7];
  assign regs$008 = regs[  8];
  assign regs$009 = regs[  9];
  assign regs$010 = regs[ 10];
  assign regs$011 = regs[ 11];
  assign regs$012 = regs[ 12];
  assign regs$013 = regs[ 13];
  assign regs$014 = regs[ 14];
  assign regs$015 = regs[ 15];
  logic   [   3:0] write_addr[0:0];
  assign write_addr[  0] = write_addr$000;
  logic   [   0:0] write_call[0:0];
  assign write_call[  0] = write_call$000;
  logic   [ 141:0] write_data[0:0];
  assign write_data[  0] = write_data$000;

  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def handle_writes():
  //         for i in range(num_write_ports):
  //           if s.write_call[i]:
  //             s.regs[s.write_addr[i]].n = s.write_data[i]

  // logic for handle_writes()
  always @ (posedge clk) begin
    for (i=0; i < num_write_ports; i=i+1)
    begin
      if (write_call[i]) begin
        regs[write_addr[i]] <= write_data[i];
      end
      else begin
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_reads():
  //         for i in range(num_read_ports):
  //           s.read_data[i].v = s.regs[s.read_addr[i]]

  // logic for handle_reads()
  always @ (*) begin
    for (i=0; i < num_read_ports; i=i+1)
    begin
      read_data[i] = regs[read_addr[i]];
    end
  end


endmodule // AsynchronousRAM_0x3c5ad87dd535d6cd

//-----------------------------------------------------------------------------
// Mux_0x71ecd1c0a6217ee5
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.mux {"dtype": 1, "nports": 16}
// PyMTL: verilator_xinit = zeros
module Mux_0x71ecd1c0a6217ee5
(
  input  logic [   0:0] clk,
  input  logic [   0:0] mux_in_$000,
  input  logic [   0:0] mux_in_$010,
  input  logic [   0:0] mux_in_$011,
  input  logic [   0:0] mux_in_$012,
  input  logic [   0:0] mux_in_$013,
  input  logic [   0:0] mux_in_$014,
  input  logic [   0:0] mux_in_$015,
  input  logic [   0:0] mux_in_$001,
  input  logic [   0:0] mux_in_$002,
  input  logic [   0:0] mux_in_$003,
  input  logic [   0:0] mux_in_$004,
  input  logic [   0:0] mux_in_$005,
  input  logic [   0:0] mux_in_$006,
  input  logic [   0:0] mux_in_$007,
  input  logic [   0:0] mux_in_$008,
  input  logic [   0:0] mux_in_$009,
  output logic  [   0:0] mux_out,
  input  logic [   3:0] mux_select,
  input  logic [   0:0] reset
);

  // localparam declarations
  localparam nports = 16;


  // array declarations
  logic   [   0:0] mux_in_[0:15];
  assign mux_in_[  0] = mux_in_$000;
  assign mux_in_[  1] = mux_in_$001;
  assign mux_in_[  2] = mux_in_$002;
  assign mux_in_[  3] = mux_in_$003;
  assign mux_in_[  4] = mux_in_$004;
  assign mux_in_[  5] = mux_in_$005;
  assign mux_in_[  6] = mux_in_$006;
  assign mux_in_[  7] = mux_in_$007;
  assign mux_in_[  8] = mux_in_$008;
  assign mux_in_[  9] = mux_in_$009;
  assign mux_in_[ 10] = mux_in_$010;
  assign mux_in_[ 11] = mux_in_$011;
  assign mux_in_[ 12] = mux_in_$012;
  assign mux_in_[ 13] = mux_in_$013;
  assign mux_in_[ 14] = mux_in_$014;
  assign mux_in_[ 15] = mux_in_$015;

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def select():
  //       assert s.mux_select < nports
  //       s.mux_out.v = s.mux_in_[s.mux_select]

  // logic for select()
  always @ (*) begin
    mux_out = mux_in_[mux_select];
  end


endmodule // Mux_0x71ecd1c0a6217ee5

//-----------------------------------------------------------------------------
// Fetch_0x4aa1acfe24534b0
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: core.rtl.frontend.fetch {"MemMsg": "MemMsg: op: 1 ts: 2 ad: 64 da: 8", "fetch_interface": "peek <R> () -> (msg: Bits(162)); take <C> () -> ()"}
// PyMTL: verilator_xinit = zeros
module Fetch_0x4aa1acfe24534b0
(
  input  logic [   0:0] check_redirect_redirect,
  input  logic [  63:0] check_redirect_target,
  input  logic [   0:0] clk,
  output logic [   0:0] mem_recv_call,
  input  logic [  75:0] mem_recv_msg,
  input  logic [   0:0] mem_recv_rdy,
  output logic [   0:0] mem_send_call,
  output logic  [ 135:0] mem_send_msg,
  input  logic [   0:0] mem_send_rdy,
  output logic [ 161:0] peek_msg,
  output logic  [   0:0] peek_rdy,
  input  logic [   0:0] reset,
  input  logic [   0:0] take_call
);

  // logic declarations
  logic   [  63:0] drop_unit_output_data_data;


  // register declarations
  logic    [   0:0] advance_f0;
  logic    [   0:0] advance_f1;
  logic    [   0:0] drop_unit$drop_call;
  logic    [   0:0] drop_unit$output_call;
  logic    [   0:0] fetch_msg$write_call;
  logic    [ 161:0] fetch_msg$write_data;
  logic    [   0:0] fetch_val$write_call;
  logic    [   0:0] fetch_val$write_data;
  logic    [  31:0] inst_from_mem;
  logic    [   0:0] pc$write_call;
  logic    [  63:0] pc$write_data;

  // localparam declarations
  localparam ACCESS_FAULT = 2'd2;
  localparam ADDRESS_MISALIGNED = 2'd1;
  localparam INSTRUCTION_ACCESS_FAULT = 4'd1;
  localparam INSTRUCTION_ADDRESS_MISALIGNED = 4'd0;
  localparam OK = 2'd0;
  localparam PIPELINE_MSG_STATUS_EXCEPTION_RAISED = 2'd1;
  localparam PIPELINE_MSG_STATUS_VALID = 2'd0;
  localparam ilen = 32;
  localparam ilen_bytes = 4;

  // fetch_val temporaries
  logic   [   0:0] fetch_val$clk;
  logic   [   0:0] fetch_val$reset;
  logic   [   0:0] fetch_val$read_data;

  Register_0x19ffe7c045ca5b3a fetch_val
  (
    .clk        ( fetch_val$clk ),
    .write_call ( fetch_val$write_call ),
    .write_data ( fetch_val$write_data ),
    .reset      ( fetch_val$reset ),
    .read_data  ( fetch_val$read_data )
  );

  // pc temporaries
  logic   [   0:0] pc$clk;
  logic   [   0:0] pc$reset;
  logic   [  63:0] pc$read_data;

  Register_0x11f1129223d5cba0 pc
  (
    .clk        ( pc$clk ),
    .write_call ( pc$write_call ),
    .write_data ( pc$write_data ),
    .reset      ( pc$reset ),
    .read_data  ( pc$read_data )
  );

  // drop_unit temporaries
  logic   [  75:0] drop_unit$input_data;
  logic   [   0:0] drop_unit$clk;
  logic   [   0:0] drop_unit$input_rdy;
  logic   [   0:0] drop_unit$reset;
  logic   [   0:0] drop_unit$output_rdy;
  logic   [   0:0] drop_unit$drop_rdy;
  logic   [   0:0] drop_unit$input_call;
  logic   [  75:0] drop_unit$output_data;
  logic   [   0:0] drop_unit$drop_status_occurred;

  DropUnit_0x1ffc4326f33abd32 drop_unit
  (
    .input_data           ( drop_unit$input_data ),
    .output_call          ( drop_unit$output_call ),
    .clk                  ( drop_unit$clk ),
    .input_rdy            ( drop_unit$input_rdy ),
    .drop_call            ( drop_unit$drop_call ),
    .reset                ( drop_unit$reset ),
    .output_rdy           ( drop_unit$output_rdy ),
    .drop_rdy             ( drop_unit$drop_rdy ),
    .input_call           ( drop_unit$input_call ),
    .output_data          ( drop_unit$output_data ),
    .drop_status_occurred ( drop_unit$drop_status_occurred )
  );

  // in_flight temporaries
  logic   [   0:0] in_flight$clk;
  logic   [   0:0] in_flight$write_call;
  logic   [   0:0] in_flight$write_data;
  logic   [   0:0] in_flight$reset;
  logic   [   0:0] in_flight$read_data;

  Register_0x19ffe7c045ca5b3a in_flight
  (
    .clk        ( in_flight$clk ),
    .write_call ( in_flight$write_call ),
    .write_data ( in_flight$write_data ),
    .reset      ( in_flight$reset ),
    .read_data  ( in_flight$read_data )
  );

  // fetch_msg temporaries
  logic   [   0:0] fetch_msg$clk;
  logic   [   0:0] fetch_msg$reset;
  logic   [ 161:0] fetch_msg$read_data;

  Register_0x538c25b0b2fe6de fetch_msg
  (
    .clk        ( fetch_msg$clk ),
    .write_call ( fetch_msg$write_call ),
    .write_data ( fetch_msg$write_data ),
    .reset      ( fetch_msg$reset ),
    .read_data  ( fetch_msg$read_data )
  );

  // signal connections
  assign drop_unit$clk              = clk;
  assign drop_unit$input_data       = mem_recv_msg;
  assign drop_unit$input_rdy        = mem_recv_rdy;
  assign drop_unit$reset            = reset;
  assign drop_unit_output_data_data = drop_unit$output_data[63:0];
  assign fetch_msg$clk              = clk;
  assign fetch_msg$reset            = reset;
  assign fetch_val$clk              = clk;
  assign fetch_val$reset            = reset;
  assign in_flight$clk              = clk;
  assign in_flight$reset            = reset;
  assign in_flight$write_call       = advance_f0;
  assign in_flight$write_data       = 1'd1;
  assign mem_recv_call              = drop_unit$input_call;
  assign mem_send_call              = advance_f0;
  assign mem_send_msg[135:132]      = 4'd0;
  assign mem_send_msg[66:64]        = 3'd4;
  assign pc$clk                     = clk;
  assign pc$reset                   = reset;
  assign peek_msg                   = fetch_msg$read_data;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def pymtl_is_broken_connect_does_not_work():
  //       s.inst_from_mem.v = s.drop_unit_output_data_data[0:ilen]

  // logic for pymtl_is_broken_connect_does_not_work()
  always @ (*) begin
    inst_from_mem = drop_unit_output_data_data[(ilen)-1:0];
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_advance():
  //       s.advance_f1.v = s.drop_unit.output_rdy and (not s.fetch_val.read_data or
  //                                                    s.take_call)
  //       s.advance_f0.v = not s.in_flight.read_data or s.drop_unit.drop_status_occurred or s.advance_f1

  // logic for handle_advance()
  always @ (*) begin
    advance_f1 = (drop_unit$output_rdy&&(!fetch_val$read_data||take_call));
    advance_f0 = (!in_flight$read_data||drop_unit$drop_status_occurred||advance_f1);
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_redirect():
  //       if s.check_redirect_redirect:
  //         # drop if in flight
  //         s.drop_unit.drop_call.v = s.in_flight.read_data
  //         # the new PC is the target
  //         s.pc.write_data.v = s.check_redirect_target
  //         s.pc.write_call.v = 1
  //
  //       else:
  //         s.drop_unit.drop_call.v = 0
  //         # if we are issuing now, the new PC is just ilen_bytes more than the last one
  //         # Insert BTB here!
  //         s.pc.write_data.v = s.pc.read_data + ilen_bytes
  //         s.pc.write_call.v = s.advance_f0

  // logic for handle_redirect()
  always @ (*) begin
    if (check_redirect_redirect) begin
      drop_unit$drop_call = in_flight$read_data;
      pc$write_data = check_redirect_target;
      pc$write_call = 1;
    end
    else begin
      drop_unit$drop_call = 0;
      pc$write_data = (pc$read_data+ilen_bytes);
      pc$write_call = advance_f0;
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_f1():
  //       s.fetch_val.write_call.v = 0
  //       s.fetch_val.write_data.v = 0
  //       s.fetch_msg.write_call.v = 0
  //       s.fetch_msg.write_data.v = 0
  //       s.drop_unit.output_call.v = 0
  //
  //       if s.check_redirect_redirect:
  //         # invalidate the output
  //         s.peek_rdy.v = 0
  //         # write a 0 into the valid register
  //         s.fetch_val.write_call.v = 1
  //       else:
  //         s.peek_rdy.v = s.fetch_val.read_data
  //
  //         if s.drop_unit.output_rdy and (not s.fetch_val.read_data or
  //                                        s.take_call):
  //           s.fetch_val.write_call.v = 1
  //           s.fetch_val.write_data.v = 1
  //           s.fetch_msg.write_call.v = 1
  //           s.drop_unit.output_call.v = 1
  //
  //           s.fetch_msg.write_data.hdr_pc.v = s.pc.read_data
  //           if s.drop_unit.output_data.stat != MemMsgStatus.OK:
  //             s.fetch_msg.write_data.hdr_status.v = PipelineMsgStatus.PIPELINE_MSG_STATUS_EXCEPTION_RAISED
  //             if s.drop_unit.output_data.stat == MemMsgStatus.ADDRESS_MISALIGNED:
  //               s.fetch_msg.write_data.exception_info_mcause.v = ExceptionCode.INSTRUCTION_ADDRESS_MISALIGNED
  //             elif s.drop_unit.output_data.stat == MemMsgStatus.ACCESS_FAULT:
  //               s.fetch_msg.write_data.exception_info_mcause.v = ExceptionCode.INSTRUCTION_ACCESS_FAULT
  //             # save the faulting PC as mtval
  //             s.fetch_msg.write_data.exception_info_mtval.v = s.pc.read_data
  //           else:
  //             s.fetch_msg.write_data.hdr_status.v = PipelineMsgStatus.PIPELINE_MSG_STATUS_VALID
  //             s.fetch_msg.write_data.inst.v = s.inst_from_mem
  //             s.fetch_msg.write_data.pc_succ.v = s.pc.write_data
  //         elif s.take_call:
  //           # someone is calling, but we are stalled, so give them output but
  //           # unset valid
  //           s.fetch_val.write_call.v = 1
  //           s.fetch_val.write_data.v = 0

  // logic for handle_f1()
  always @ (*) begin
    fetch_val$write_call = 0;
    fetch_val$write_data = 0;
    fetch_msg$write_call = 0;
    fetch_msg$write_data = 0;
    drop_unit$output_call = 0;
    if (check_redirect_redirect) begin
      peek_rdy = 0;
      fetch_val$write_call = 1;
    end
    else begin
      peek_rdy = fetch_val$read_data;
      if ((drop_unit$output_rdy&&(!fetch_val$read_data||take_call))) begin
        fetch_val$write_call = 1;
        fetch_val$write_data = 1;
        fetch_msg$write_call = 1;
        drop_unit$output_call = 1;
        fetch_msg$write_data[(66)-1:2] = pc$read_data;
        if ((drop_unit$output_data[(69)-1:67] != OK)) begin
          fetch_msg$write_data[(2)-1:0] = PIPELINE_MSG_STATUS_EXCEPTION_RAISED;
          if ((drop_unit$output_data[(69)-1:67] == ADDRESS_MISALIGNED)) begin
            fetch_msg$write_data[(70)-1:66] = INSTRUCTION_ADDRESS_MISALIGNED;
          end
          else begin
            if ((drop_unit$output_data[(69)-1:67] == ACCESS_FAULT)) begin
              fetch_msg$write_data[(70)-1:66] = INSTRUCTION_ACCESS_FAULT;
            end
            else begin
            end
          end
          fetch_msg$write_data[(134)-1:70] = pc$read_data;
        end
        else begin
          fetch_msg$write_data[(2)-1:0] = PIPELINE_MSG_STATUS_VALID;
          fetch_msg$write_data[(98)-1:66] = inst_from_mem;
          fetch_msg$write_data[(162)-1:98] = pc$write_data;
        end
      end
      else begin
        if (take_call) begin
          fetch_val$write_call = 1;
          fetch_val$write_data = 0;
        end
        else begin
        end
      end
    end
  end

  // PYMTL SOURCE:
  //
  // @s.combinational
  // def write_addr():
  //       s.mem_send_msg.addr.v = s.pc.write_data

  // logic for write_addr()
  always @ (*) begin
    mem_send_msg[(131)-1:67] = pc$write_data;
  end


endmodule // Fetch_0x4aa1acfe24534b0

//-----------------------------------------------------------------------------
// Register_0x11f1129223d5cba0
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(64)); write <C> (data: Bits(64)) -> ()", "reset_value": 0}
// PyMTL: verilator_xinit = zeros
module Register_0x11f1129223d5cba0
(
  input  logic [   0:0] clk,
  output logic [  63:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [  63:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [  63:0] reg_value;

  // localparam declarations
  localparam reset_value = 0;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.reset:
  //           s.reg_value.n = reset_value
  //         elif s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (reset) begin
      reg_value <= reset_value;
    end
    else begin
      if (update) begin
        reg_value <= write_data;
      end
      else begin
      end
    end
  end


endmodule // Register_0x11f1129223d5cba0

//-----------------------------------------------------------------------------
// DropUnit_0x1ffc4326f33abd32
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.drop_unit {"interface": "drop <CR> () -> (); drop_status () -> (occurred: Bits(1)); output <CR> () -> (data: Bits(76))"}
// PyMTL: verilator_xinit = zeros
module DropUnit_0x1ffc4326f33abd32
(
  input  logic [   0:0] clk,
  input  logic [   0:0] drop_call,
  output logic  [   0:0] drop_rdy,
  output logic  [   0:0] drop_status_occurred,
  output logic  [   0:0] input_call,
  input  logic [  75:0] input_data,
  input  logic [   0:0] input_rdy,
  input  logic [   0:0] output_call,
  output logic [  75:0] output_data,
  output logic  [   0:0] output_rdy,
  input  logic [   0:0] reset
);

  // register declarations
  logic    [   0:0] drop_pending$write_data;
  logic    [   0:0] drop_pending_curr;

  // drop_pending temporaries
  logic   [   0:0] drop_pending$clk;
  logic   [   0:0] drop_pending$reset;
  logic   [   0:0] drop_pending$read_data;

  Register_0x360ff20b8ea9d7d7 drop_pending
  (
    .clk        ( drop_pending$clk ),
    .write_data ( drop_pending$write_data ),
    .reset      ( drop_pending$reset ),
    .read_data  ( drop_pending$read_data )
  );

  // signal connections
  assign drop_pending$clk   = clk;
  assign drop_pending$reset = reset;
  assign output_data        = input_data;


  // PYMTL SOURCE:
  //
  // @s.combinational
  // def handle_drop():
  //       s.drop_pending_curr.v = s.drop_pending.read_data or s.drop_call
  //       s.drop_status_occurred.v = s.drop_pending_curr and s.input_rdy
  //       s.drop_rdy.v = not s.drop_pending.read_data
  //
  //       if s.drop_status_occurred:
  //         s.input_call.v = 1
  //         s.output_rdy.v = 0
  //         s.drop_pending.write_data.v = 0
  //       elif s.drop_pending_curr:
  //         s.input_call.v = 0
  //         s.output_rdy.v = 0
  //         s.drop_pending.write_data.v = 1
  //       else:
  //         s.input_call.v = s.output_call
  //         s.output_rdy.v = s.input_rdy
  //         s.drop_pending.write_data.v = 0

  // logic for handle_drop()
  always @ (*) begin
    drop_pending_curr = (drop_pending$read_data||drop_call);
    drop_status_occurred = (drop_pending_curr&&input_rdy);
    drop_rdy = !drop_pending$read_data;
    if (drop_status_occurred) begin
      input_call = 1;
      output_rdy = 0;
      drop_pending$write_data = 0;
    end
    else begin
      if (drop_pending_curr) begin
        input_call = 0;
        output_rdy = 0;
        drop_pending$write_data = 1;
      end
      else begin
        input_call = output_call;
        output_rdy = input_rdy;
        drop_pending$write_data = 0;
      end
    end
  end


endmodule // DropUnit_0x1ffc4326f33abd32

//-----------------------------------------------------------------------------
// Register_0x538c25b0b2fe6de
//-----------------------------------------------------------------------------
// PyMTL: dump_vcd = False
// PyMTL: util.rtl.register {"interface": "read () -> (data: Bits(162)); write <C> (data: Bits(162)) -> ()", "reset_value": null}
// PyMTL: verilator_xinit = zeros
module Register_0x538c25b0b2fe6de
(
  input  logic [   0:0] clk,
  output logic [ 161:0] read_data,
  input  logic [   0:0] reset,
  input  logic [   0:0] write_call,
  input  logic [ 161:0] write_data
);

  // logic declarations
  logic   [   0:0] update;


  // register declarations
  logic    [ 161:0] reg_value;

  // signal connections
  assign read_data = reg_value;
  assign update    = write_call;


  // PYMTL SOURCE:
  //
  // @s.tick_rtl
  // def update():
  //         if s.update:
  //           s.reg_value.n = s.write_data

  // logic for update()
  always @ (posedge clk) begin
    if (update) begin
      reg_value <= write_data;
    end
    else begin
    end
  end


endmodule // Register_0x538c25b0b2fe6de

